`timescale 1ns / 10ps

module tt_um_gray_sobel (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire LFSR_enable_i_sync;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire net142;
 wire _0043_;
 wire net143;
 wire _0045_;
 wire net144;
 wire _0047_;
 wire net145;
 wire _0049_;
 wire net146;
 wire _0051_;
 wire net147;
 wire _0053_;
 wire _0054_;
 wire net148;
 wire _0056_;
 wire net149;
 wire _0058_;
 wire net150;
 wire _0060_;
 wire net151;
 wire _0062_;
 wire net152;
 wire _0064_;
 wire net153;
 wire _0066_;
 wire net154;
 wire _0068_;
 wire net155;
 wire _0070_;
 wire net156;
 wire _0072_;
 wire net157;
 wire _0074_;
 wire net158;
 wire _0076_;
 wire net159;
 wire _0078_;
 wire net160;
 wire _0080_;
 wire net161;
 wire _0082_;
 wire net162;
 wire _0084_;
 wire net163;
 wire _0086_;
 wire net164;
 wire _0088_;
 wire net165;
 wire _0090_;
 wire net166;
 wire _0092_;
 wire net167;
 wire _0094_;
 wire net168;
 wire _0096_;
 wire net169;
 wire _0098_;
 wire net170;
 wire _0100_;
 wire clknet_leaf_0_clk;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire net138;
 wire frame_done_i_sync;
 wire \gray_sobel0.gray_scale0.nreset_i ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[0] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[1] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[2] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[3] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[4] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[5] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[6] ;
 wire \gray_sobel0.gray_scale0.out_px_gray_o[7] ;
 wire \gray_sobel0.gray_scale0.px_rdy_i ;
 wire \gray_sobel0.gray_scale0.px_rdy_o ;
 wire \gray_sobel0.out_px_sobel[0] ;
 wire \gray_sobel0.out_px_sobel[1] ;
 wire \gray_sobel0.out_px_sobel[2] ;
 wire \gray_sobel0.out_px_sobel[3] ;
 wire \gray_sobel0.out_px_sobel[4] ;
 wire \gray_sobel0.out_px_sobel[5] ;
 wire \gray_sobel0.out_px_sobel[6] ;
 wire \gray_sobel0.out_px_sobel[7] ;
 wire \gray_sobel0.px_rdy_o_sobel ;
 wire \gray_sobel0.select_sobel_mux ;
 wire \gray_sobel0.sobel0.counter_pixels[0] ;
 wire \gray_sobel0.sobel0.counter_pixels[10] ;
 wire \gray_sobel0.sobel0.counter_pixels[11] ;
 wire \gray_sobel0.sobel0.counter_pixels[12] ;
 wire \gray_sobel0.sobel0.counter_pixels[13] ;
 wire \gray_sobel0.sobel0.counter_pixels[14] ;
 wire \gray_sobel0.sobel0.counter_pixels[15] ;
 wire \gray_sobel0.sobel0.counter_pixels[16] ;
 wire \gray_sobel0.sobel0.counter_pixels[17] ;
 wire \gray_sobel0.sobel0.counter_pixels[18] ;
 wire \gray_sobel0.sobel0.counter_pixels[19] ;
 wire \gray_sobel0.sobel0.counter_pixels[1] ;
 wire \gray_sobel0.sobel0.counter_pixels[20] ;
 wire \gray_sobel0.sobel0.counter_pixels[21] ;
 wire \gray_sobel0.sobel0.counter_pixels[22] ;
 wire \gray_sobel0.sobel0.counter_pixels[23] ;
 wire \gray_sobel0.sobel0.counter_pixels[2] ;
 wire \gray_sobel0.sobel0.counter_pixels[3] ;
 wire \gray_sobel0.sobel0.counter_pixels[4] ;
 wire \gray_sobel0.sobel0.counter_pixels[5] ;
 wire \gray_sobel0.sobel0.counter_pixels[6] ;
 wire \gray_sobel0.sobel0.counter_pixels[7] ;
 wire \gray_sobel0.sobel0.counter_pixels[8] ;
 wire \gray_sobel0.sobel0.counter_pixels[9] ;
 wire \gray_sobel0.sobel0.counter_sobel[0] ;
 wire \gray_sobel0.sobel0.counter_sobel[1] ;
 wire \gray_sobel0.sobel0.counter_sobel[2] ;
 wire \gray_sobel0.sobel0.counter_sobel[3] ;
 wire \gray_sobel0.sobel0.fsm_state[0] ;
 wire \gray_sobel0.sobel0.fsm_state[1] ;
 wire \gray_sobel0.sobel0.next[0] ;
 wire \gray_sobel0.sobel0.next[1] ;
 wire \gray_sobel0.sobel0.px_ready ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i0[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i1[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i2[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i3[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i4[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i5[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i7[7] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[5] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ;
 wire \gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ;
 wire in_data_rdy;
 wire in_lfsr_rdy;
 wire \input_data[0] ;
 wire \input_data[10] ;
 wire \input_data[11] ;
 wire \input_data[12] ;
 wire \input_data[13] ;
 wire \input_data[14] ;
 wire \input_data[15] ;
 wire \input_data[16] ;
 wire \input_data[17] ;
 wire \input_data[18] ;
 wire \input_data[19] ;
 wire \input_data[1] ;
 wire \input_data[20] ;
 wire \input_data[21] ;
 wire \input_data[22] ;
 wire \input_data[23] ;
 wire \input_data[2] ;
 wire \input_data[3] ;
 wire \input_data[4] ;
 wire \input_data[5] ;
 wire \input_data[6] ;
 wire \input_data[7] ;
 wire \input_data[8] ;
 wire \input_data[9] ;
 wire \lfsr0.config_done_o ;
 wire \lfsr0.config_i ;
 wire \lfsr0.lfsr_done ;
 wire \lfsr0.lfsr_en_i ;
 wire \lfsr0.lfsr_out[0] ;
 wire \lfsr0.lfsr_out[10] ;
 wire \lfsr0.lfsr_out[11] ;
 wire \lfsr0.lfsr_out[12] ;
 wire \lfsr0.lfsr_out[13] ;
 wire \lfsr0.lfsr_out[14] ;
 wire \lfsr0.lfsr_out[15] ;
 wire \lfsr0.lfsr_out[16] ;
 wire \lfsr0.lfsr_out[17] ;
 wire \lfsr0.lfsr_out[18] ;
 wire \lfsr0.lfsr_out[19] ;
 wire \lfsr0.lfsr_out[1] ;
 wire \lfsr0.lfsr_out[20] ;
 wire \lfsr0.lfsr_out[21] ;
 wire \lfsr0.lfsr_out[22] ;
 wire \lfsr0.lfsr_out[23] ;
 wire \lfsr0.lfsr_out[2] ;
 wire \lfsr0.lfsr_out[3] ;
 wire \lfsr0.lfsr_out[4] ;
 wire \lfsr0.lfsr_out[5] ;
 wire \lfsr0.lfsr_out[6] ;
 wire \lfsr0.lfsr_out[7] ;
 wire \lfsr0.lfsr_out[8] ;
 wire \lfsr0.lfsr_out[9] ;
 wire \lfsr0.lfsr_rdy_o ;
 wire \lfsr0.seed_reg[0] ;
 wire \lfsr0.seed_reg[10] ;
 wire \lfsr0.seed_reg[11] ;
 wire \lfsr0.seed_reg[12] ;
 wire \lfsr0.seed_reg[13] ;
 wire \lfsr0.seed_reg[14] ;
 wire \lfsr0.seed_reg[15] ;
 wire \lfsr0.seed_reg[16] ;
 wire \lfsr0.seed_reg[17] ;
 wire \lfsr0.seed_reg[18] ;
 wire \lfsr0.seed_reg[19] ;
 wire \lfsr0.seed_reg[1] ;
 wire \lfsr0.seed_reg[20] ;
 wire \lfsr0.seed_reg[21] ;
 wire \lfsr0.seed_reg[22] ;
 wire \lfsr0.seed_reg[23] ;
 wire \lfsr0.seed_reg[2] ;
 wire \lfsr0.seed_reg[3] ;
 wire \lfsr0.seed_reg[4] ;
 wire \lfsr0.seed_reg[5] ;
 wire \lfsr0.seed_reg[6] ;
 wire \lfsr0.seed_reg[7] ;
 wire \lfsr0.seed_reg[8] ;
 wire \lfsr0.seed_reg[9] ;
 wire \lfsr0.stop_reg[0] ;
 wire \lfsr0.stop_reg[10] ;
 wire \lfsr0.stop_reg[11] ;
 wire \lfsr0.stop_reg[12] ;
 wire \lfsr0.stop_reg[13] ;
 wire \lfsr0.stop_reg[14] ;
 wire \lfsr0.stop_reg[15] ;
 wire \lfsr0.stop_reg[16] ;
 wire \lfsr0.stop_reg[17] ;
 wire \lfsr0.stop_reg[18] ;
 wire \lfsr0.stop_reg[19] ;
 wire \lfsr0.stop_reg[1] ;
 wire \lfsr0.stop_reg[20] ;
 wire \lfsr0.stop_reg[21] ;
 wire \lfsr0.stop_reg[22] ;
 wire \lfsr0.stop_reg[23] ;
 wire \lfsr0.stop_reg[2] ;
 wire \lfsr0.stop_reg[3] ;
 wire \lfsr0.stop_reg[4] ;
 wire \lfsr0.stop_reg[5] ;
 wire \lfsr0.stop_reg[6] ;
 wire \lfsr0.stop_reg[7] ;
 wire \lfsr0.stop_reg[8] ;
 wire \lfsr0.stop_reg[9] ;
 wire lfsr_mode_sel_i_sync;
 wire \nreset_sync0.r_sync ;
 wire \sa0.clear_i ;
 wire \sa0.en_i ;
 wire \sa0.signature_o[0] ;
 wire \sa0.signature_o[10] ;
 wire \sa0.signature_o[11] ;
 wire \sa0.signature_o[12] ;
 wire \sa0.signature_o[13] ;
 wire \sa0.signature_o[14] ;
 wire \sa0.signature_o[15] ;
 wire \sa0.signature_o[16] ;
 wire \sa0.signature_o[17] ;
 wire \sa0.signature_o[18] ;
 wire \sa0.signature_o[19] ;
 wire \sa0.signature_o[1] ;
 wire \sa0.signature_o[20] ;
 wire \sa0.signature_o[21] ;
 wire \sa0.signature_o[22] ;
 wire \sa0.signature_o[23] ;
 wire \sa0.signature_o[2] ;
 wire \sa0.signature_o[3] ;
 wire \sa0.signature_o[4] ;
 wire \sa0.signature_o[5] ;
 wire \sa0.signature_o[6] ;
 wire \sa0.signature_o[7] ;
 wire \sa0.signature_o[8] ;
 wire \sa0.signature_o[9] ;
 wire \sgnl_sync0.signal_sync ;
 wire \sgnl_sync1.signal_o ;
 wire \sgnl_sync1.signal_sync ;
 wire \sgnl_sync2.signal_sync ;
 wire \sgnl_sync3.signal_sync ;
 wire \sgnl_sync4.signal_sync ;
 wire \sgnl_sync5.signal_sync ;
 wire \sgnl_sync6.signal_sync ;
 wire \sgnl_sync7.signal_sync ;
 wire \sgnl_sync8.signal_sync ;
 wire \spi0.data_tx[0] ;
 wire \spi0.data_tx[10] ;
 wire \spi0.data_tx[11] ;
 wire \spi0.data_tx[12] ;
 wire \spi0.data_tx[13] ;
 wire \spi0.data_tx[14] ;
 wire \spi0.data_tx[15] ;
 wire \spi0.data_tx[16] ;
 wire \spi0.data_tx[17] ;
 wire \spi0.data_tx[18] ;
 wire \spi0.data_tx[19] ;
 wire \spi0.data_tx[1] ;
 wire \spi0.data_tx[20] ;
 wire \spi0.data_tx[21] ;
 wire \spi0.data_tx[22] ;
 wire \spi0.data_tx[23] ;
 wire \spi0.data_tx[2] ;
 wire \spi0.data_tx[3] ;
 wire \spi0.data_tx[4] ;
 wire \spi0.data_tx[5] ;
 wire \spi0.data_tx[6] ;
 wire \spi0.data_tx[7] ;
 wire \spi0.data_tx[8] ;
 wire \spi0.data_tx[9] ;
 wire \spi0.rxtx_done ;
 wire \spi0.rxtx_done_reg ;
 wire \spi0.rxtx_done_rising ;
 wire \spi0.signal_sync1.async_signal_i ;
 wire \spi0.signal_sync1.signal_sync ;
 wire \spi0.spi0.counter[0] ;
 wire \spi0.spi0.counter[1] ;
 wire \spi0.spi0.counter[2] ;
 wire \spi0.spi0.counter[3] ;
 wire \spi0.spi0.counter[4] ;
 wire \spi0.spi0.counter[5] ;
 wire \spi0.spi0.data_rx_o[0] ;
 wire \spi0.spi0.data_rx_o[10] ;
 wire \spi0.spi0.data_rx_o[11] ;
 wire \spi0.spi0.data_rx_o[12] ;
 wire \spi0.spi0.data_rx_o[13] ;
 wire \spi0.spi0.data_rx_o[14] ;
 wire \spi0.spi0.data_rx_o[15] ;
 wire \spi0.spi0.data_rx_o[16] ;
 wire \spi0.spi0.data_rx_o[17] ;
 wire \spi0.spi0.data_rx_o[18] ;
 wire \spi0.spi0.data_rx_o[19] ;
 wire \spi0.spi0.data_rx_o[1] ;
 wire \spi0.spi0.data_rx_o[20] ;
 wire \spi0.spi0.data_rx_o[21] ;
 wire \spi0.spi0.data_rx_o[22] ;
 wire \spi0.spi0.data_rx_o[23] ;
 wire \spi0.spi0.data_rx_o[2] ;
 wire \spi0.spi0.data_rx_o[3] ;
 wire \spi0.spi0.data_rx_o[4] ;
 wire \spi0.spi0.data_rx_o[5] ;
 wire \spi0.spi0.data_rx_o[6] ;
 wire \spi0.spi0.data_rx_o[7] ;
 wire \spi0.spi0.data_rx_o[8] ;
 wire \spi0.spi0.data_rx_o[9] ;
 wire \spi0.spi0.sdo_o ;
 wire \spi0.spi0.sdo_register[0] ;
 wire \spi0.spi0.sdo_register[10] ;
 wire \spi0.spi0.sdo_register[11] ;
 wire \spi0.spi0.sdo_register[12] ;
 wire \spi0.spi0.sdo_register[13] ;
 wire \spi0.spi0.sdo_register[14] ;
 wire \spi0.spi0.sdo_register[15] ;
 wire \spi0.spi0.sdo_register[16] ;
 wire \spi0.spi0.sdo_register[17] ;
 wire \spi0.spi0.sdo_register[18] ;
 wire \spi0.spi0.sdo_register[19] ;
 wire \spi0.spi0.sdo_register[1] ;
 wire \spi0.spi0.sdo_register[20] ;
 wire \spi0.spi0.sdo_register[21] ;
 wire \spi0.spi0.sdo_register[22] ;
 wire \spi0.spi0.sdo_register[2] ;
 wire \spi0.spi0.sdo_register[3] ;
 wire \spi0.spi0.sdo_register[4] ;
 wire \spi0.spi0.sdo_register[5] ;
 wire \spi0.spi0.sdo_register[6] ;
 wire \spi0.spi0.sdo_register[7] ;
 wire \spi0.spi0.sdo_register[8] ;
 wire \spi0.spi0.sdo_register[9] ;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net139;
 wire net140;
 wire net141;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire [1:0] clknet_0_ui_in;
 wire [1:0] clknet_2_0__leaf_ui_in;
 wire [1:0] clknet_2_1__leaf_ui_in;
 wire [1:0] clknet_2_2__leaf_ui_in;
 wire [1:0] clknet_2_3__leaf_ui_in;

 sky130_fd_sc_hd__inv_2 _1348_ (.A(net123),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1349_ (.A(\gray_sobel0.sobel0.fsm_state[1] ),
    .Y(_1140_));
 sky130_fd_sc_hd__inv_2 _1350_ (.A(net74),
    .Y(_1141_));
 sky130_fd_sc_hd__inv_2 _1351_ (.A(\lfsr0.stop_reg[0] ),
    .Y(_1142_));
 sky130_fd_sc_hd__inv_2 _1352_ (.A(\lfsr0.lfsr_out[0] ),
    .Y(_1143_));
 sky130_fd_sc_hd__inv_2 _1353_ (.A(\lfsr0.lfsr_out[3] ),
    .Y(_1144_));
 sky130_fd_sc_hd__inv_2 _1354_ (.A(\lfsr0.lfsr_out[5] ),
    .Y(_1145_));
 sky130_fd_sc_hd__inv_2 _1355_ (.A(\lfsr0.stop_reg[6] ),
    .Y(_1146_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(\lfsr0.stop_reg[7] ),
    .Y(_1147_));
 sky130_fd_sc_hd__inv_2 _1357_ (.A(\lfsr0.lfsr_out[9] ),
    .Y(_1148_));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(\lfsr0.lfsr_out[10] ),
    .Y(_1149_));
 sky130_fd_sc_hd__inv_2 _1359_ (.A(\lfsr0.lfsr_out[11] ),
    .Y(_1150_));
 sky130_fd_sc_hd__inv_2 _1360_ (.A(\lfsr0.lfsr_out[14] ),
    .Y(_1151_));
 sky130_fd_sc_hd__inv_2 _1361_ (.A(\lfsr0.lfsr_out[15] ),
    .Y(_1152_));
 sky130_fd_sc_hd__inv_2 _1362_ (.A(\lfsr0.lfsr_out[16] ),
    .Y(_1153_));
 sky130_fd_sc_hd__inv_2 _1363_ (.A(\lfsr0.stop_reg[17] ),
    .Y(_1154_));
 sky130_fd_sc_hd__inv_2 _1364_ (.A(\lfsr0.stop_reg[20] ),
    .Y(_1155_));
 sky130_fd_sc_hd__inv_2 _1365_ (.A(\lfsr0.stop_reg[23] ),
    .Y(_1156_));
 sky130_fd_sc_hd__inv_2 _1366_ (.A(net68),
    .Y(_1157_));
 sky130_fd_sc_hd__inv_2 _1367_ (.A(net276),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1368_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[5] ),
    .Y(_1158_));
 sky130_fd_sc_hd__inv_2 _1369_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ),
    .Y(_1159_));
 sky130_fd_sc_hd__inv_2 _1370_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[5] ),
    .Y(_1160_));
 sky130_fd_sc_hd__inv_2 _1371_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[2] ),
    .Y(_1161_));
 sky130_fd_sc_hd__inv_2 _1372_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[6] ),
    .Y(_1162_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[5] ),
    .Y(_1163_));
 sky130_fd_sc_hd__inv_2 _1374_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[4] ),
    .Y(_1164_));
 sky130_fd_sc_hd__inv_2 _1375_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[3] ),
    .Y(_1165_));
 sky130_fd_sc_hd__inv_2 _2647__2 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _1377_ (.A(\gray_sobel0.sobel0.px_ready ),
    .Y(_1166_));
 sky130_fd_sc_hd__or4_1 _1378_ (.A(\gray_sobel0.sobel0.counter_pixels[5] ),
    .B(\gray_sobel0.sobel0.counter_pixels[4] ),
    .C(\gray_sobel0.sobel0.counter_pixels[7] ),
    .D(\gray_sobel0.sobel0.counter_pixels[6] ),
    .X(_1167_));
 sky130_fd_sc_hd__or4b_1 _1379_ (.A(\gray_sobel0.sobel0.counter_pixels[1] ),
    .B(\gray_sobel0.sobel0.counter_pixels[3] ),
    .C(\gray_sobel0.sobel0.counter_pixels[2] ),
    .D_N(\gray_sobel0.sobel0.counter_pixels[0] ),
    .X(_1168_));
 sky130_fd_sc_hd__or4_1 _1380_ (.A(\gray_sobel0.sobel0.counter_pixels[13] ),
    .B(\gray_sobel0.sobel0.counter_pixels[12] ),
    .C(\gray_sobel0.sobel0.counter_pixels[15] ),
    .D(\gray_sobel0.sobel0.counter_pixels[14] ),
    .X(_1169_));
 sky130_fd_sc_hd__or4_1 _1381_ (.A(\gray_sobel0.sobel0.counter_pixels[9] ),
    .B(\gray_sobel0.sobel0.counter_pixels[8] ),
    .C(\gray_sobel0.sobel0.counter_pixels[11] ),
    .D(\gray_sobel0.sobel0.counter_pixels[10] ),
    .X(_1170_));
 sky130_fd_sc_hd__or4_1 _1382_ (.A(\gray_sobel0.sobel0.counter_pixels[17] ),
    .B(\gray_sobel0.sobel0.counter_pixels[16] ),
    .C(\gray_sobel0.sobel0.counter_pixels[19] ),
    .D(\gray_sobel0.sobel0.counter_pixels[18] ),
    .X(_1171_));
 sky130_fd_sc_hd__or4_1 _1383_ (.A(\gray_sobel0.sobel0.counter_pixels[21] ),
    .B(\gray_sobel0.sobel0.counter_pixels[20] ),
    .C(\gray_sobel0.sobel0.counter_pixels[23] ),
    .D(\gray_sobel0.sobel0.counter_pixels[22] ),
    .X(_1172_));
 sky130_fd_sc_hd__or3_1 _1384_ (.A(_1169_),
    .B(_1170_),
    .C(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__nor4_1 _1385_ (.A(_1167_),
    .B(_1168_),
    .C(_1171_),
    .D(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nor2_1 _1386_ (.A(\gray_sobel0.sobel0.fsm_state[1] ),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__or2_1 _1387_ (.A(\gray_sobel0.sobel0.fsm_state[1] ),
    .B(net197),
    .X(_1176_));
 sky130_fd_sc_hd__a21oi_1 _1388_ (.A1(\gray_sobel0.sobel0.fsm_state[1] ),
    .A2(net197),
    .B1(\gray_sobel0.sobel0.fsm_state[0] ),
    .Y(_1177_));
 sky130_fd_sc_hd__a22o_2 _1389_ (.A1(\gray_sobel0.sobel0.fsm_state[0] ),
    .A2(_1175_),
    .B1(_1176_),
    .B2(_1177_),
    .X(\gray_sobel0.sobel0.next[0] ));
 sky130_fd_sc_hd__and3b_1 _1390_ (.A_N(\gray_sobel0.sobel0.fsm_state[0] ),
    .B(\gray_sobel0.sobel0.fsm_state[1] ),
    .C(net6),
    .X(_1178_));
 sky130_fd_sc_hd__a31o_1 _1391_ (.A1(\gray_sobel0.sobel0.fsm_state[0] ),
    .A2(_1140_),
    .A3(_1174_),
    .B1(_1178_),
    .X(\gray_sobel0.sobel0.next[1] ));
 sky130_fd_sc_hd__and2_1 _1392_ (.A(net440),
    .B(net74),
    .X(in_lfsr_rdy));
 sky130_fd_sc_hd__mux2_1 _1393_ (.A0(in_data_rdy),
    .A1(net282),
    .S(net74),
    .X(\gray_sobel0.gray_scale0.px_rdy_i ));
 sky130_fd_sc_hd__a2bb2o_1 _1394_ (.A1_N(_1147_),
    .A2_N(\lfsr0.lfsr_out[7] ),
    .B1(\lfsr0.stop_reg[14] ),
    .B2(_1151_),
    .X(_1179_));
 sky130_fd_sc_hd__o22a_1 _1395_ (.A1(\lfsr0.stop_reg[5] ),
    .A2(_1145_),
    .B1(\lfsr0.stop_reg[14] ),
    .B2(_1151_),
    .X(_1180_));
 sky130_fd_sc_hd__xor2_1 _1396_ (.A(\lfsr0.stop_reg[22] ),
    .B(\lfsr0.lfsr_out[22] ),
    .X(_1181_));
 sky130_fd_sc_hd__xnor2_1 _1397_ (.A(\lfsr0.stop_reg[12] ),
    .B(\lfsr0.lfsr_out[12] ),
    .Y(_1182_));
 sky130_fd_sc_hd__xor2_1 _1398_ (.A(\lfsr0.stop_reg[4] ),
    .B(\lfsr0.lfsr_out[4] ),
    .X(_1183_));
 sky130_fd_sc_hd__xnor2_1 _1399_ (.A(\lfsr0.stop_reg[2] ),
    .B(\lfsr0.lfsr_out[2] ),
    .Y(_1184_));
 sky130_fd_sc_hd__nand2_1 _1400_ (.A(\lfsr0.stop_reg[1] ),
    .B(\lfsr0.lfsr_out[1] ),
    .Y(_1185_));
 sky130_fd_sc_hd__or2_1 _1401_ (.A(\lfsr0.stop_reg[1] ),
    .B(\lfsr0.lfsr_out[1] ),
    .X(_1186_));
 sky130_fd_sc_hd__or2_1 _1402_ (.A(\lfsr0.stop_reg[21] ),
    .B(\lfsr0.lfsr_out[21] ),
    .X(_1187_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(\lfsr0.stop_reg[21] ),
    .B(\lfsr0.lfsr_out[21] ),
    .Y(_1188_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(\lfsr0.stop_reg[13] ),
    .B(\lfsr0.lfsr_out[13] ),
    .Y(_1189_));
 sky130_fd_sc_hd__or2_1 _1405_ (.A(\lfsr0.stop_reg[13] ),
    .B(\lfsr0.lfsr_out[13] ),
    .X(_1190_));
 sky130_fd_sc_hd__a221o_1 _1406_ (.A1(_1187_),
    .A2(_1188_),
    .B1(_1189_),
    .B2(_1190_),
    .C1(_1181_),
    .X(_1191_));
 sky130_fd_sc_hd__a221o_1 _1407_ (.A1(\lfsr0.stop_reg[10] ),
    .A2(_1149_),
    .B1(_1185_),
    .B2(_1186_),
    .C1(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__a22o_1 _1408_ (.A1(_1146_),
    .A2(\lfsr0.lfsr_out[6] ),
    .B1(_1156_),
    .B2(\lfsr0.lfsr_out[23] ),
    .X(_1193_));
 sky130_fd_sc_hd__a221o_1 _1409_ (.A1(\lfsr0.stop_reg[5] ),
    .A2(_1145_),
    .B1(_1147_),
    .B2(\lfsr0.lfsr_out[7] ),
    .C1(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__a2bb2o_1 _1410_ (.A1_N(\lfsr0.stop_reg[9] ),
    .A2_N(_1148_),
    .B1(\lfsr0.stop_reg[11] ),
    .B2(_1150_),
    .X(_1195_));
 sky130_fd_sc_hd__a221o_1 _1411_ (.A1(_1142_),
    .A2(\lfsr0.lfsr_out[0] ),
    .B1(\lfsr0.stop_reg[16] ),
    .B2(_1153_),
    .C1(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__xor2_1 _1412_ (.A(\lfsr0.stop_reg[19] ),
    .B(\lfsr0.lfsr_out[19] ),
    .X(_1197_));
 sky130_fd_sc_hd__a221o_1 _1413_ (.A1(\lfsr0.stop_reg[0] ),
    .A2(_1143_),
    .B1(\lfsr0.stop_reg[15] ),
    .B2(_1152_),
    .C1(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__xor2_1 _1414_ (.A(\lfsr0.stop_reg[18] ),
    .B(\lfsr0.lfsr_out[18] ),
    .X(_1199_));
 sky130_fd_sc_hd__xor2_1 _1415_ (.A(\lfsr0.stop_reg[8] ),
    .B(\lfsr0.lfsr_out[8] ),
    .X(_1200_));
 sky130_fd_sc_hd__or4_1 _1416_ (.A(_1196_),
    .B(_1198_),
    .C(_1199_),
    .D(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__a2bb2o_1 _1417_ (.A1_N(\lfsr0.lfsr_out[6] ),
    .A2_N(_1146_),
    .B1(_1144_),
    .B2(\lfsr0.stop_reg[3] ),
    .X(_1202_));
 sky130_fd_sc_hd__a221o_1 _1418_ (.A1(_1154_),
    .A2(\lfsr0.lfsr_out[17] ),
    .B1(_1155_),
    .B2(\lfsr0.lfsr_out[20] ),
    .C1(_1179_),
    .X(_1203_));
 sky130_fd_sc_hd__a2111o_1 _1419_ (.A1(\lfsr0.stop_reg[9] ),
    .A2(_1148_),
    .B1(_1183_),
    .C1(_1202_),
    .D1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__o221a_1 _1420_ (.A1(\lfsr0.stop_reg[3] ),
    .A2(_1144_),
    .B1(\lfsr0.stop_reg[16] ),
    .B2(_1153_),
    .C1(_1182_),
    .X(_1205_));
 sky130_fd_sc_hd__o211a_1 _1421_ (.A1(\lfsr0.stop_reg[11] ),
    .A2(_1150_),
    .B1(_1180_),
    .C1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__o221a_1 _1422_ (.A1(\lfsr0.stop_reg[15] ),
    .A2(_1152_),
    .B1(_1156_),
    .B2(\lfsr0.lfsr_out[23] ),
    .C1(_1184_),
    .X(_1207_));
 sky130_fd_sc_hd__o22a_1 _1423_ (.A1(\lfsr0.stop_reg[10] ),
    .A2(_1149_),
    .B1(_1155_),
    .B2(\lfsr0.lfsr_out[20] ),
    .X(_1208_));
 sky130_fd_sc_hd__o211a_1 _1424_ (.A1(_1154_),
    .A2(\lfsr0.lfsr_out[17] ),
    .B1(_1207_),
    .C1(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__and3b_1 _1425_ (.A_N(_1204_),
    .B(_1206_),
    .C(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__or4b_1 _1426_ (.A(_1192_),
    .B(_1194_),
    .C(_1201_),
    .D_N(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__inv_2 _1427_ (.A(net32),
    .Y(\lfsr0.lfsr_done ));
 sky130_fd_sc_hd__nor2_1 _1428_ (.A(_1157_),
    .B(\lfsr0.lfsr_done ),
    .Y(_0000_));
 sky130_fd_sc_hd__or3b_1 _1429_ (.A(\spi0.spi0.counter[2] ),
    .B(\spi0.spi0.counter[5] ),
    .C_N(\spi0.spi0.counter[3] ),
    .X(_1212_));
 sky130_fd_sc_hd__and4bb_1 _1430_ (.A_N(\spi0.spi0.counter[1] ),
    .B_N(_1212_),
    .C(_0002_),
    .D(\spi0.spi0.counter[4] ),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _1431_ (.A(\spi0.data_tx[16] ),
    .B(net50),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(net273),
    .A1(\spi0.data_tx[17] ),
    .S(net50),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1433_ (.A0(net257),
    .A1(\spi0.data_tx[18] ),
    .S(net50),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(net266),
    .A1(\spi0.data_tx[19] ),
    .S(net50),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1435_ (.A0(net262),
    .A1(\spi0.data_tx[20] ),
    .S(net50),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1436_ (.A0(net261),
    .A1(\spi0.data_tx[21] ),
    .S(net50),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1437_ (.A0(net268),
    .A1(\spi0.data_tx[22] ),
    .S(net53),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(net258),
    .A1(\spi0.data_tx[23] ),
    .S(net50),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(net252),
    .A1(\spi0.data_tx[8] ),
    .S(net53),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(net255),
    .A1(\spi0.data_tx[9] ),
    .S(net52),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(net263),
    .A1(\spi0.data_tx[10] ),
    .S(net51),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(net269),
    .A1(\spi0.data_tx[11] ),
    .S(net51),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _1443_ (.A0(net256),
    .A1(\spi0.data_tx[12] ),
    .S(net51),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(net271),
    .A1(\spi0.data_tx[13] ),
    .S(net51),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(net259),
    .A1(\spi0.data_tx[14] ),
    .S(net51),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _1446_ (.A0(net272),
    .A1(\spi0.data_tx[15] ),
    .S(net51),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _1447_ (.A0(net253),
    .A1(\spi0.data_tx[0] ),
    .S(net51),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _1448_ (.A0(net251),
    .A1(\spi0.data_tx[1] ),
    .S(net51),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _1449_ (.A0(net264),
    .A1(\spi0.data_tx[2] ),
    .S(net51),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _1450_ (.A0(net254),
    .A1(\spi0.data_tx[3] ),
    .S(net51),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(net270),
    .A1(\spi0.data_tx[4] ),
    .S(net52),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(net260),
    .A1(\spi0.data_tx[5] ),
    .S(net52),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1453_ (.A0(net265),
    .A1(\spi0.data_tx[6] ),
    .S(net52),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1454_ (.A0(net250),
    .A1(\spi0.data_tx[7] ),
    .S(net52),
    .X(_0024_));
 sky130_fd_sc_hd__xor2_1 _1455_ (.A(net305),
    .B(net276),
    .X(_0003_));
 sky130_fd_sc_hd__and3_1 _1456_ (.A(\spi0.spi0.counter[1] ),
    .B(\spi0.spi0.counter[0] ),
    .C(\spi0.spi0.counter[2] ),
    .X(_1213_));
 sky130_fd_sc_hd__a21oi_1 _1457_ (.A1(\spi0.spi0.counter[1] ),
    .A2(\spi0.spi0.counter[0] ),
    .B1(net289),
    .Y(_1214_));
 sky130_fd_sc_hd__nor2_1 _1458_ (.A(_1213_),
    .B(net290),
    .Y(_0004_));
 sky130_fd_sc_hd__and2_1 _1459_ (.A(\spi0.spi0.counter[3] ),
    .B(_1213_),
    .X(_1215_));
 sky130_fd_sc_hd__nor2_1 _1460_ (.A(net50),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__o21a_1 _1461_ (.A1(net278),
    .A2(_1213_),
    .B1(_1216_),
    .X(_0005_));
 sky130_fd_sc_hd__or2_1 _1462_ (.A(\spi0.spi0.counter[4] ),
    .B(_1215_),
    .X(_1217_));
 sky130_fd_sc_hd__nand2_1 _1463_ (.A(\spi0.spi0.counter[4] ),
    .B(_1215_),
    .Y(_1218_));
 sky130_fd_sc_hd__and3b_1 _1464_ (.A_N(net50),
    .B(_1217_),
    .C(_1218_),
    .X(_0006_));
 sky130_fd_sc_hd__xnor2_1 _1465_ (.A(net275),
    .B(_1218_),
    .Y(_0007_));
 sky130_fd_sc_hd__and2b_1 _1466_ (.A_N(\spi0.rxtx_done_reg ),
    .B(\spi0.rxtx_done ),
    .X(\spi0.rxtx_done_rising ));
 sky130_fd_sc_hd__nor2_1 _1467_ (.A(net33),
    .B(net47),
    .Y(_1219_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(\gray_sobel0.gray_scale0.px_rdy_o ),
    .A1(\gray_sobel0.gray_scale0.px_rdy_i ),
    .S(net77),
    .X(_1220_));
 sky130_fd_sc_hd__and2b_1 _1469_ (.A_N(\sgnl_sync1.signal_o ),
    .B(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__o21ai_4 _1470_ (.A1(net33),
    .A2(net47),
    .B1(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__or4b_2 _1471_ (.A(\gray_sobel0.sobel0.counter_sobel[0] ),
    .B(\gray_sobel0.sobel0.counter_sobel[2] ),
    .C(\gray_sobel0.sobel0.counter_sobel[3] ),
    .D_N(\gray_sobel0.sobel0.counter_sobel[1] ),
    .X(_1223_));
 sky130_fd_sc_hd__or2_1 _1472_ (.A(\gray_sobel0.sobel0.counter_sobel[1] ),
    .B(\gray_sobel0.sobel0.counter_sobel[0] ),
    .X(_1224_));
 sky130_fd_sc_hd__or3b_1 _1473_ (.A(_1224_),
    .B(\gray_sobel0.sobel0.counter_sobel[2] ),
    .C_N(\gray_sobel0.sobel0.counter_sobel[3] ),
    .X(_1225_));
 sky130_fd_sc_hd__a22o_1 _1474_ (.A1(net47),
    .A2(_1223_),
    .B1(_1225_),
    .B2(net33),
    .X(_1226_));
 sky130_fd_sc_hd__nor2_1 _1475_ (.A(_1222_),
    .B(_1226_),
    .Y(_0001_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(\input_data[4] ),
    .A1(\lfsr0.lfsr_out[4] ),
    .S(net73),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_2 _1477_ (.A0(\input_data[5] ),
    .A1(\lfsr0.lfsr_out[5] ),
    .S(net73),
    .X(_1228_));
 sky130_fd_sc_hd__and2_1 _1478_ (.A(_1227_),
    .B(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__nor2_1 _1479_ (.A(_1227_),
    .B(_1228_),
    .Y(_1230_));
 sky130_fd_sc_hd__nor2_1 _1480_ (.A(_1229_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__mux2_2 _1481_ (.A0(\input_data[9] ),
    .A1(\lfsr0.lfsr_out[9] ),
    .S(net73),
    .X(_1232_));
 sky130_fd_sc_hd__xnor2_1 _1482_ (.A(_1231_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(\input_data[12] ),
    .A1(\lfsr0.lfsr_out[12] ),
    .S(net72),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(\input_data[18] ),
    .A1(\lfsr0.lfsr_out[18] ),
    .S(net74),
    .X(_1235_));
 sky130_fd_sc_hd__nor2_1 _1485_ (.A(_1234_),
    .B(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__and2_1 _1486_ (.A(_1234_),
    .B(_1235_),
    .X(_1237_));
 sky130_fd_sc_hd__nor2_1 _1487_ (.A(_1236_),
    .B(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__mux2_2 _1488_ (.A0(\input_data[21] ),
    .A1(\lfsr0.lfsr_out[21] ),
    .S(net72),
    .X(_1239_));
 sky130_fd_sc_hd__xor2_1 _1489_ (.A(_1238_),
    .B(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__and2b_1 _1490_ (.A_N(_1233_),
    .B(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__xnor2_1 _1491_ (.A(_1233_),
    .B(_1240_),
    .Y(_0033_));
 sky130_fd_sc_hd__mux2_2 _1492_ (.A0(\input_data[6] ),
    .A1(\lfsr0.lfsr_out[6] ),
    .S(net73),
    .X(_1242_));
 sky130_fd_sc_hd__nand2_1 _1493_ (.A(_1228_),
    .B(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__or2_1 _1494_ (.A(_1228_),
    .B(_1242_),
    .X(_1244_));
 sky130_fd_sc_hd__nand2_1 _1495_ (.A(_1243_),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__mux2_1 _1496_ (.A0(\input_data[10] ),
    .A1(\lfsr0.lfsr_out[10] ),
    .S(net72),
    .X(_1246_));
 sky130_fd_sc_hd__xor2_1 _1497_ (.A(_1245_),
    .B(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__a21oi_1 _1498_ (.A1(_1231_),
    .A2(_1232_),
    .B1(_1229_),
    .Y(_1248_));
 sky130_fd_sc_hd__nor2_1 _1499_ (.A(_1247_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _1500_ (.A(_1247_),
    .B(_1248_),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2b_1 _1501_ (.A_N(_1249_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__mux2_2 _1502_ (.A0(\input_data[13] ),
    .A1(\lfsr0.lfsr_out[13] ),
    .S(net72),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(\input_data[19] ),
    .A1(\lfsr0.lfsr_out[19] ),
    .S(net75),
    .X(_1253_));
 sky130_fd_sc_hd__and2_1 _1504_ (.A(_1252_),
    .B(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__nor2_1 _1505_ (.A(_1252_),
    .B(_1253_),
    .Y(_1255_));
 sky130_fd_sc_hd__nor2_1 _1506_ (.A(_1254_),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__mux2_2 _1507_ (.A0(\input_data[22] ),
    .A1(\lfsr0.lfsr_out[22] ),
    .S(net72),
    .X(_1257_));
 sky130_fd_sc_hd__xor2_1 _1508_ (.A(_1256_),
    .B(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__xnor2_1 _1509_ (.A(_1251_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_1 _1510_ (.A(_1241_),
    .B(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__or2_1 _1511_ (.A(_1241_),
    .B(_1259_),
    .X(_1261_));
 sky130_fd_sc_hd__nand2_1 _1512_ (.A(_1260_),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__a21o_1 _1513_ (.A1(_1238_),
    .A2(_1239_),
    .B1(_1237_),
    .X(_1263_));
 sky130_fd_sc_hd__nand2b_1 _1514_ (.A_N(_1262_),
    .B(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__xnor2_1 _1515_ (.A(_1262_),
    .B(_1263_),
    .Y(_0034_));
 sky130_fd_sc_hd__a21o_1 _1516_ (.A1(_1256_),
    .A2(_1257_),
    .B1(_1254_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _1517_ (.A0(\input_data[14] ),
    .A1(\lfsr0.lfsr_out[14] ),
    .S(net72),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(\input_data[20] ),
    .A1(\lfsr0.lfsr_out[20] ),
    .S(net75),
    .X(_1267_));
 sky130_fd_sc_hd__nor2_1 _1519_ (.A(_1266_),
    .B(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__and2_1 _1520_ (.A(_1266_),
    .B(_1267_),
    .X(_1269_));
 sky130_fd_sc_hd__nor2_1 _1521_ (.A(_1268_),
    .B(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__mux2_2 _1522_ (.A0(\input_data[23] ),
    .A1(\lfsr0.lfsr_out[23] ),
    .S(net73),
    .X(_1271_));
 sky130_fd_sc_hd__xor2_1 _1523_ (.A(_1270_),
    .B(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_2 _1524_ (.A0(\input_data[7] ),
    .A1(\lfsr0.lfsr_out[7] ),
    .S(net73),
    .X(_1273_));
 sky130_fd_sc_hd__nand2_1 _1525_ (.A(_1242_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__or2_1 _1526_ (.A(_1242_),
    .B(_1273_),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _1527_ (.A0(\input_data[11] ),
    .A1(\lfsr0.lfsr_out[11] ),
    .S(net72),
    .X(_1276_));
 sky130_fd_sc_hd__nand3_1 _1528_ (.A(_1274_),
    .B(_1275_),
    .C(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__a21o_1 _1529_ (.A1(_1274_),
    .A2(_1275_),
    .B1(_1276_),
    .X(_1278_));
 sky130_fd_sc_hd__nand2_1 _1530_ (.A(_1277_),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__a21boi_1 _1531_ (.A1(_1244_),
    .A2(_1246_),
    .B1_N(_1243_),
    .Y(_1280_));
 sky130_fd_sc_hd__or2_1 _1532_ (.A(_1279_),
    .B(_1280_),
    .X(_1281_));
 sky130_fd_sc_hd__nand2_1 _1533_ (.A(_1279_),
    .B(_1280_),
    .Y(_1282_));
 sky130_fd_sc_hd__and2_1 _1534_ (.A(_1281_),
    .B(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__nand2_1 _1535_ (.A(_1272_),
    .B(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__or2_1 _1536_ (.A(_1272_),
    .B(_1283_),
    .X(_1285_));
 sky130_fd_sc_hd__nand2_1 _1537_ (.A(_1284_),
    .B(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__a21oi_1 _1538_ (.A1(_1250_),
    .A2(_1258_),
    .B1(_1249_),
    .Y(_1287_));
 sky130_fd_sc_hd__or2_1 _1539_ (.A(_1286_),
    .B(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__nand2_1 _1540_ (.A(_1286_),
    .B(_1287_),
    .Y(_1289_));
 sky130_fd_sc_hd__nand2_1 _1541_ (.A(_1288_),
    .B(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__nand2b_1 _1542_ (.A_N(_1290_),
    .B(_1265_),
    .Y(_1291_));
 sky130_fd_sc_hd__xor2_1 _1543_ (.A(_1265_),
    .B(_1290_),
    .X(_1292_));
 sky130_fd_sc_hd__a21oi_1 _1544_ (.A1(_1260_),
    .A2(_1264_),
    .B1(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__nor2_1 _1545_ (.A(_1234_),
    .B(_1273_),
    .Y(_1294_));
 sky130_fd_sc_hd__and2_1 _1546_ (.A(_1234_),
    .B(_1273_),
    .X(_1295_));
 sky130_fd_sc_hd__nor2_1 _1547_ (.A(_1294_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__mux2_2 _1548_ (.A0(\input_data[15] ),
    .A1(\lfsr0.lfsr_out[15] ),
    .S(net72),
    .X(_1297_));
 sky130_fd_sc_hd__xnor2_1 _1549_ (.A(_1296_),
    .B(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__a21o_1 _1550_ (.A1(_1274_),
    .A2(_1277_),
    .B1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__nand3_1 _1551_ (.A(_1274_),
    .B(_1277_),
    .C(_1298_),
    .Y(_1300_));
 sky130_fd_sc_hd__and2_1 _1552_ (.A(_1299_),
    .B(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__or2_1 _1553_ (.A(_1239_),
    .B(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__nand2_1 _1554_ (.A(_1239_),
    .B(_1301_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2_1 _1555_ (.A(_1302_),
    .B(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__a21oi_1 _1556_ (.A1(_1281_),
    .A2(_1284_),
    .B1(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__and3_1 _1557_ (.A(_1281_),
    .B(_1284_),
    .C(_1304_),
    .X(_1306_));
 sky130_fd_sc_hd__or2_1 _1558_ (.A(_1305_),
    .B(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__a21o_1 _1559_ (.A1(_1270_),
    .A2(_1271_),
    .B1(_1269_),
    .X(_1308_));
 sky130_fd_sc_hd__and2b_1 _1560_ (.A_N(_1307_),
    .B(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__xor2_1 _1561_ (.A(_1307_),
    .B(_1308_),
    .X(_1310_));
 sky130_fd_sc_hd__a21oi_1 _1562_ (.A1(_1288_),
    .A2(_1291_),
    .B1(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__and3_1 _1563_ (.A(_1288_),
    .B(_1291_),
    .C(_1310_),
    .X(_1312_));
 sky130_fd_sc_hd__or2_1 _1564_ (.A(_1311_),
    .B(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__nor3b_1 _1565_ (.A(_1311_),
    .B(_1312_),
    .C_N(_1293_),
    .Y(_1314_));
 sky130_fd_sc_hd__xnor2_1 _1566_ (.A(_1293_),
    .B(_1313_),
    .Y(_0036_));
 sky130_fd_sc_hd__xnor2_1 _1567_ (.A(_1252_),
    .B(_1257_),
    .Y(_1315_));
 sky130_fd_sc_hd__a21oi_1 _1568_ (.A1(_1296_),
    .A2(_1297_),
    .B1(_1295_),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2_1 _1569_ (.A(_1315_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__or2_1 _1570_ (.A(_1315_),
    .B(_1316_),
    .X(_1318_));
 sky130_fd_sc_hd__nand2_1 _1571_ (.A(_1317_),
    .B(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__a21oi_1 _1572_ (.A1(_1299_),
    .A2(_1303_),
    .B1(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__and3_1 _1573_ (.A(_1299_),
    .B(_1303_),
    .C(_1319_),
    .X(_1321_));
 sky130_fd_sc_hd__nor2_1 _1574_ (.A(_1320_),
    .B(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__o21a_1 _1575_ (.A1(_1305_),
    .A2(_1309_),
    .B1(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__nor3_1 _1576_ (.A(_1305_),
    .B(_1309_),
    .C(_1322_),
    .Y(_1324_));
 sky130_fd_sc_hd__nor2_1 _1577_ (.A(_1323_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__o21a_1 _1578_ (.A1(_1311_),
    .A2(_1314_),
    .B1(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__nor3_1 _1579_ (.A(_1311_),
    .B(_1314_),
    .C(_1325_),
    .Y(_1327_));
 sky130_fd_sc_hd__nor2_1 _1580_ (.A(_1326_),
    .B(_1327_),
    .Y(_0037_));
 sky130_fd_sc_hd__nor2_1 _1581_ (.A(_1266_),
    .B(_1271_),
    .Y(_1328_));
 sky130_fd_sc_hd__and2_1 _1582_ (.A(_1266_),
    .B(_1271_),
    .X(_1329_));
 sky130_fd_sc_hd__and4bb_1 _1583_ (.A_N(_1328_),
    .B_N(_1329_),
    .C(_1252_),
    .D(_1257_),
    .X(_1330_));
 sky130_fd_sc_hd__o2bb2a_1 _1584_ (.A1_N(_1252_),
    .A2_N(_1257_),
    .B1(_1328_),
    .B2(_1329_),
    .X(_1331_));
 sky130_fd_sc_hd__nor2_1 _1585_ (.A(_1330_),
    .B(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__and2b_1 _1586_ (.A_N(_1318_),
    .B(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__nand2_1 _1587_ (.A(_1320_),
    .B(_1332_),
    .Y(_1334_));
 sky130_fd_sc_hd__or2_1 _1588_ (.A(_1320_),
    .B(_1332_),
    .X(_1335_));
 sky130_fd_sc_hd__nand2_1 _1589_ (.A(_1334_),
    .B(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hd__a21oi_1 _1590_ (.A1(_1318_),
    .A2(_1336_),
    .B1(_1333_),
    .Y(_1337_));
 sky130_fd_sc_hd__o21ai_1 _1591_ (.A1(_1323_),
    .A2(_1326_),
    .B1(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__or3_1 _1592_ (.A(_1323_),
    .B(_1326_),
    .C(_1337_),
    .X(_1339_));
 sky130_fd_sc_hd__and2_1 _1593_ (.A(_1338_),
    .B(_1339_),
    .X(_0038_));
 sky130_fd_sc_hd__o21a_1 _1594_ (.A1(_1329_),
    .A2(_1330_),
    .B1(_1297_),
    .X(_1340_));
 sky130_fd_sc_hd__nor3_1 _1595_ (.A(_1297_),
    .B(_1329_),
    .C(_1330_),
    .Y(_1341_));
 sky130_fd_sc_hd__nor2_1 _1596_ (.A(_1340_),
    .B(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__xnor2_1 _1597_ (.A(_1333_),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__a21oi_1 _1598_ (.A1(_1334_),
    .A2(_1338_),
    .B1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__and3_1 _1599_ (.A(_1334_),
    .B(_1338_),
    .C(_1343_),
    .X(_1345_));
 sky130_fd_sc_hd__nor2_1 _1600_ (.A(_1344_),
    .B(_1345_),
    .Y(_0039_));
 sky130_fd_sc_hd__a211o_1 _1601_ (.A1(_1333_),
    .A2(_1342_),
    .B1(_1344_),
    .C1(_1340_),
    .X(_0040_));
 sky130_fd_sc_hd__and3_1 _1602_ (.A(_1260_),
    .B(_1264_),
    .C(_1292_),
    .X(_1346_));
 sky130_fd_sc_hd__nor2_1 _1603_ (.A(_1293_),
    .B(_1346_),
    .Y(_0035_));
 sky130_fd_sc_hd__mux2_1 _1604_ (.A0(\input_data[0] ),
    .A1(\spi0.spi0.data_rx_o[16] ),
    .S(net65),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1605_ (.A0(net434),
    .A1(\spi0.spi0.data_rx_o[17] ),
    .S(net65),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(net428),
    .A1(\spi0.spi0.data_rx_o[18] ),
    .S(net63),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(net411),
    .A1(\spi0.spi0.data_rx_o[19] ),
    .S(net63),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(net394),
    .A1(\spi0.spi0.data_rx_o[20] ),
    .S(net65),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(net441),
    .A1(\spi0.spi0.data_rx_o[21] ),
    .S(net64),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(net458),
    .A1(\spi0.spi0.data_rx_o[22] ),
    .S(net64),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1611_ (.A0(\input_data[7] ),
    .A1(\spi0.spi0.data_rx_o[23] ),
    .S(net65),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1612_ (.A0(\input_data[8] ),
    .A1(\spi0.spi0.data_rx_o[8] ),
    .S(net64),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1613_ (.A0(\input_data[9] ),
    .A1(\spi0.spi0.data_rx_o[9] ),
    .S(net64),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(\input_data[10] ),
    .A1(\spi0.spi0.data_rx_o[10] ),
    .S(net63),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _1615_ (.A0(\input_data[11] ),
    .A1(\spi0.spi0.data_rx_o[11] ),
    .S(net63),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(\input_data[12] ),
    .A1(\spi0.spi0.data_rx_o[12] ),
    .S(net63),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _1617_ (.A0(net423),
    .A1(\spi0.spi0.data_rx_o[13] ),
    .S(net63),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _1618_ (.A0(net433),
    .A1(\spi0.spi0.data_rx_o[14] ),
    .S(net63),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _1619_ (.A0(\input_data[15] ),
    .A1(\spi0.spi0.data_rx_o[15] ),
    .S(net63),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _1620_ (.A0(net412),
    .A1(\spi0.spi0.data_rx_o[0] ),
    .S(net65),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _1621_ (.A0(net442),
    .A1(\spi0.spi0.data_rx_o[1] ),
    .S(net64),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(net437),
    .A1(\spi0.spi0.data_rx_o[2] ),
    .S(net64),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(net432),
    .A1(\spi0.spi0.data_rx_o[3] ),
    .S(net64),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _1624_ (.A0(net429),
    .A1(\spi0.spi0.data_rx_o[4] ),
    .S(net64),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _1625_ (.A0(net444),
    .A1(\spi0.spi0.data_rx_o[5] ),
    .S(net63),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _1626_ (.A0(net452),
    .A1(\spi0.spi0.data_rx_o[6] ),
    .S(net63),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _1627_ (.A0(net449),
    .A1(\spi0.spi0.data_rx_o[7] ),
    .S(net64),
    .X(_0149_));
 sky130_fd_sc_hd__and4bb_1 _1628_ (.A_N(net74),
    .B_N(lfsr_mode_sel_i_sync),
    .C(frame_done_i_sync),
    .D(\sa0.en_i ),
    .X(_0378_));
 sky130_fd_sc_hd__and4b_1 _1629_ (.A_N(lfsr_mode_sel_i_sync),
    .B(\lfsr0.lfsr_done ),
    .C(net74),
    .D(\sa0.en_i ),
    .X(_0379_));
 sky130_fd_sc_hd__a21o_1 _1630_ (.A1(_1157_),
    .A2(_0379_),
    .B1(_0378_),
    .X(_0380_));
 sky130_fd_sc_hd__a21oi_1 _1631_ (.A1(_1141_),
    .A2(lfsr_mode_sel_i_sync),
    .B1(\sa0.en_i ),
    .Y(_0381_));
 sky130_fd_sc_hd__o21a_2 _1632_ (.A1(_1141_),
    .A2(lfsr_mode_sel_i_sync),
    .B1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _1633_ (.A0(\gray_sobel0.px_rdy_o_sobel ),
    .A1(_1220_),
    .S(\sgnl_sync1.signal_o ),
    .X(_0383_));
 sky130_fd_sc_hd__nor3b_1 _1634_ (.A(\sa0.en_i ),
    .B(lfsr_mode_sel_i_sync),
    .C_N(net75),
    .Y(_0384_));
 sky130_fd_sc_hd__a221o_1 _1635_ (.A1(_0382_),
    .A2(_0383_),
    .B1(net62),
    .B2(\lfsr0.config_done_o ),
    .C1(_0378_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_1 _1636_ (.A(_0379_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__or2_1 _1637_ (.A(_0379_),
    .B(_0385_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _1638_ (.A0(\lfsr0.seed_reg[0] ),
    .A1(\lfsr0.stop_reg[0] ),
    .S(net70),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _1639_ (.A0(\input_data[0] ),
    .A1(\lfsr0.lfsr_out[0] ),
    .S(net73),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_2 _1640_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[0] ),
    .A1(_0389_),
    .S(net77),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _1641_ (.A0(\gray_sobel0.out_px_sobel[0] ),
    .A1(_0390_),
    .S(net76),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _1642_ (.A1(net61),
    .A2(_0388_),
    .B1(_0391_),
    .B2(_0382_),
    .X(_0392_));
 sky130_fd_sc_hd__a211o_1 _1643_ (.A1(\sa0.signature_o[0] ),
    .A2(net22),
    .B1(net19),
    .C1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__o21a_1 _1644_ (.A1(net307),
    .A2(net15),
    .B1(_0393_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _1645_ (.A0(\lfsr0.seed_reg[1] ),
    .A1(\lfsr0.stop_reg[1] ),
    .S(net70),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _1646_ (.A0(\input_data[1] ),
    .A1(\lfsr0.lfsr_out[1] ),
    .S(net72),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_2 _1647_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[1] ),
    .A1(_0395_),
    .S(net77),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _1648_ (.A0(\gray_sobel0.out_px_sobel[1] ),
    .A1(_0396_),
    .S(net76),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _1649_ (.A1(net61),
    .A2(_0394_),
    .B1(_0397_),
    .B2(_0382_),
    .X(_0398_));
 sky130_fd_sc_hd__a211o_1 _1650_ (.A1(\sa0.signature_o[1] ),
    .A2(net22),
    .B1(net19),
    .C1(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__o21a_1 _1651_ (.A1(net310),
    .A2(net15),
    .B1(_0399_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(\lfsr0.seed_reg[2] ),
    .A1(\lfsr0.stop_reg[2] ),
    .S(net70),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _1653_ (.A0(\input_data[2] ),
    .A1(\lfsr0.lfsr_out[2] ),
    .S(net73),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_2 _1654_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[2] ),
    .A1(_0401_),
    .S(net77),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _1655_ (.A0(\gray_sobel0.out_px_sobel[2] ),
    .A1(_0402_),
    .S(net76),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _1656_ (.A1(net61),
    .A2(_0400_),
    .B1(_0403_),
    .B2(_0382_),
    .X(_0404_));
 sky130_fd_sc_hd__a211o_1 _1657_ (.A1(\sa0.signature_o[2] ),
    .A2(net22),
    .B1(net19),
    .C1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__o21a_1 _1658_ (.A1(net302),
    .A2(net15),
    .B1(_0405_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _1659_ (.A0(\lfsr0.seed_reg[3] ),
    .A1(\lfsr0.stop_reg[3] ),
    .S(net70),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _1660_ (.A0(\input_data[3] ),
    .A1(\lfsr0.lfsr_out[3] ),
    .S(net72),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_2 _1661_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[3] ),
    .A1(_0407_),
    .S(net77),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _1662_ (.A0(\gray_sobel0.out_px_sobel[3] ),
    .A1(_0408_),
    .S(net76),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _1663_ (.A1(net61),
    .A2(_0406_),
    .B1(_0409_),
    .B2(_0382_),
    .X(_0410_));
 sky130_fd_sc_hd__a211o_1 _1664_ (.A1(\sa0.signature_o[3] ),
    .A2(net22),
    .B1(net19),
    .C1(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__o21a_1 _1665_ (.A1(net309),
    .A2(net15),
    .B1(_0411_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _1666_ (.A0(\lfsr0.seed_reg[4] ),
    .A1(\lfsr0.stop_reg[4] ),
    .S(net70),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_2 _1667_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[4] ),
    .A1(_1227_),
    .S(net77),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(\gray_sobel0.out_px_sobel[4] ),
    .A1(_0413_),
    .S(net76),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _1669_ (.A1(net62),
    .A2(_0412_),
    .B1(_0414_),
    .B2(_0382_),
    .X(_0415_));
 sky130_fd_sc_hd__a211o_1 _1670_ (.A1(\sa0.signature_o[4] ),
    .A2(net22),
    .B1(net19),
    .C1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__o21a_1 _1671_ (.A1(net311),
    .A2(net15),
    .B1(_0416_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _1672_ (.A0(\lfsr0.seed_reg[5] ),
    .A1(\lfsr0.stop_reg[5] ),
    .S(net70),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_2 _1673_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[5] ),
    .A1(_1228_),
    .S(net77),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(\gray_sobel0.out_px_sobel[5] ),
    .A1(_0418_),
    .S(net76),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _1675_ (.A1(net61),
    .A2(_0417_),
    .B1(_0419_),
    .B2(_0382_),
    .X(_0420_));
 sky130_fd_sc_hd__a211o_1 _1676_ (.A1(\sa0.signature_o[5] ),
    .A2(net22),
    .B1(net19),
    .C1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__o21a_1 _1677_ (.A1(net303),
    .A2(net15),
    .B1(_0421_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _1678_ (.A0(\lfsr0.seed_reg[6] ),
    .A1(\lfsr0.stop_reg[6] ),
    .S(net71),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_2 _1679_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[6] ),
    .A1(_1242_),
    .S(net77),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(\gray_sobel0.out_px_sobel[6] ),
    .A1(_0423_),
    .S(net76),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _1681_ (.A1(net61),
    .A2(_0422_),
    .B1(_0424_),
    .B2(_0382_),
    .X(_0425_));
 sky130_fd_sc_hd__a211o_1 _1682_ (.A1(\sa0.signature_o[6] ),
    .A2(net22),
    .B1(net19),
    .C1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o21a_1 _1683_ (.A1(net308),
    .A2(net15),
    .B1(_0426_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(\lfsr0.seed_reg[7] ),
    .A1(\lfsr0.stop_reg[7] ),
    .S(net71),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_2 _1685_ (.A0(\gray_sobel0.gray_scale0.out_px_gray_o[7] ),
    .A1(_1273_),
    .S(net77),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(\gray_sobel0.out_px_sobel[7] ),
    .A1(_0428_),
    .S(net76),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _1687_ (.A1(net62),
    .A2(_0427_),
    .B1(_0429_),
    .B2(_0382_),
    .X(_0430_));
 sky130_fd_sc_hd__a211o_1 _1688_ (.A1(\sa0.signature_o[7] ),
    .A2(net22),
    .B1(net19),
    .C1(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__o21a_1 _1689_ (.A1(net294),
    .A2(net15),
    .B1(_0431_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1690_ (.A0(\lfsr0.seed_reg[8] ),
    .A1(\lfsr0.stop_reg[8] ),
    .S(net71),
    .X(_0432_));
 sky130_fd_sc_hd__and3_1 _1691_ (.A(net76),
    .B(net77),
    .C(_0382_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1692_ (.A0(\input_data[8] ),
    .A1(\lfsr0.lfsr_out[8] ),
    .S(net73),
    .X(_0434_));
 sky130_fd_sc_hd__a22o_1 _1693_ (.A1(net61),
    .A2(_0432_),
    .B1(net40),
    .B2(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__a211o_1 _1694_ (.A1(\sa0.signature_o[8] ),
    .A2(net20),
    .B1(net18),
    .C1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__o21a_1 _1695_ (.A1(net295),
    .A2(net14),
    .B1(_0436_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(\lfsr0.seed_reg[9] ),
    .A1(\lfsr0.stop_reg[9] ),
    .S(net69),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _1697_ (.A1(_1232_),
    .A2(net41),
    .B1(_0437_),
    .B2(net60),
    .X(_0438_));
 sky130_fd_sc_hd__a211o_1 _1698_ (.A1(\sa0.signature_o[9] ),
    .A2(net20),
    .B1(net18),
    .C1(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__o21a_1 _1699_ (.A1(net316),
    .A2(net14),
    .B1(_0439_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _1700_ (.A0(\lfsr0.seed_reg[10] ),
    .A1(\lfsr0.stop_reg[10] ),
    .S(net69),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _1701_ (.A1(_1246_),
    .A2(net40),
    .B1(_0440_),
    .B2(net60),
    .X(_0441_));
 sky130_fd_sc_hd__a211o_1 _1702_ (.A1(\sa0.signature_o[10] ),
    .A2(net20),
    .B1(net17),
    .C1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__o21a_1 _1703_ (.A1(net306),
    .A2(net15),
    .B1(_0442_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(\lfsr0.seed_reg[11] ),
    .A1(\lfsr0.stop_reg[11] ),
    .S(net70),
    .X(_0443_));
 sky130_fd_sc_hd__a22o_1 _1705_ (.A1(_1276_),
    .A2(net40),
    .B1(_0443_),
    .B2(net60),
    .X(_0444_));
 sky130_fd_sc_hd__a211o_1 _1706_ (.A1(\sa0.signature_o[11] ),
    .A2(_0380_),
    .B1(_0386_),
    .C1(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__o21a_1 _1707_ (.A1(net312),
    .A2(net15),
    .B1(_0445_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _1708_ (.A0(\lfsr0.seed_reg[12] ),
    .A1(\lfsr0.stop_reg[12] ),
    .S(net69),
    .X(_0446_));
 sky130_fd_sc_hd__a22o_1 _1709_ (.A1(_1234_),
    .A2(net40),
    .B1(_0446_),
    .B2(net60),
    .X(_0447_));
 sky130_fd_sc_hd__a211o_1 _1710_ (.A1(\sa0.signature_o[12] ),
    .A2(net21),
    .B1(net18),
    .C1(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__o21a_1 _1711_ (.A1(net304),
    .A2(net16),
    .B1(_0448_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _1712_ (.A0(\lfsr0.seed_reg[13] ),
    .A1(\lfsr0.stop_reg[13] ),
    .S(net69),
    .X(_0449_));
 sky130_fd_sc_hd__a22o_1 _1713_ (.A1(_1252_),
    .A2(net40),
    .B1(_0449_),
    .B2(net60),
    .X(_0450_));
 sky130_fd_sc_hd__a211o_1 _1714_ (.A1(\sa0.signature_o[13] ),
    .A2(net21),
    .B1(net17),
    .C1(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__o21a_1 _1715_ (.A1(net298),
    .A2(net14),
    .B1(_0451_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _1716_ (.A0(\lfsr0.seed_reg[14] ),
    .A1(\lfsr0.stop_reg[14] ),
    .S(net69),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _1717_ (.A1(_1266_),
    .A2(net40),
    .B1(_0452_),
    .B2(net60),
    .X(_0453_));
 sky130_fd_sc_hd__a211o_1 _1718_ (.A1(\sa0.signature_o[14] ),
    .A2(net20),
    .B1(net18),
    .C1(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__o21a_1 _1719_ (.A1(net334),
    .A2(net16),
    .B1(_0454_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(\lfsr0.seed_reg[15] ),
    .A1(\lfsr0.stop_reg[15] ),
    .S(net69),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _1721_ (.A1(_1297_),
    .A2(net40),
    .B1(_0455_),
    .B2(net60),
    .X(_0456_));
 sky130_fd_sc_hd__a211o_1 _1722_ (.A1(\sa0.signature_o[15] ),
    .A2(net20),
    .B1(net18),
    .C1(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__o21a_1 _1723_ (.A1(net299),
    .A2(net14),
    .B1(_0457_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _1724_ (.A0(\input_data[16] ),
    .A1(\lfsr0.lfsr_out[16] ),
    .S(net74),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _1725_ (.A0(\lfsr0.seed_reg[16] ),
    .A1(\lfsr0.stop_reg[16] ),
    .S(net71),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _1726_ (.A1(net41),
    .A2(_0458_),
    .B1(_0459_),
    .B2(net61),
    .X(_0460_));
 sky130_fd_sc_hd__a211o_1 _1727_ (.A1(\sa0.signature_o[16] ),
    .A2(net20),
    .B1(net17),
    .C1(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__o21a_1 _1728_ (.A1(net280),
    .A2(net16),
    .B1(_0461_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _1729_ (.A(\sa0.signature_o[17] ),
    .B(net21),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _1730_ (.A0(\input_data[17] ),
    .A1(\lfsr0.lfsr_out[17] ),
    .S(net74),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _1731_ (.A0(\lfsr0.seed_reg[17] ),
    .A1(\lfsr0.stop_reg[17] ),
    .S(net71),
    .X(_0464_));
 sky130_fd_sc_hd__a221o_1 _1732_ (.A1(net41),
    .A2(_0463_),
    .B1(_0464_),
    .B2(net62),
    .C1(net17),
    .X(_0465_));
 sky130_fd_sc_hd__o22a_1 _1733_ (.A1(net287),
    .A2(net14),
    .B1(_0462_),
    .B2(_0465_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _1734_ (.A0(\lfsr0.seed_reg[18] ),
    .A1(\lfsr0.stop_reg[18] ),
    .S(net71),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _1735_ (.A1(_1235_),
    .A2(net41),
    .B1(_0466_),
    .B2(net61),
    .X(_0467_));
 sky130_fd_sc_hd__a211o_1 _1736_ (.A1(\sa0.signature_o[18] ),
    .A2(net21),
    .B1(net17),
    .C1(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__o21a_1 _1737_ (.A1(net335),
    .A2(net14),
    .B1(_0468_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _1738_ (.A0(\lfsr0.seed_reg[19] ),
    .A1(\lfsr0.stop_reg[19] ),
    .S(net71),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _1739_ (.A1(_1253_),
    .A2(net41),
    .B1(_0469_),
    .B2(net61),
    .X(_0470_));
 sky130_fd_sc_hd__a211o_1 _1740_ (.A1(\sa0.signature_o[19] ),
    .A2(net21),
    .B1(net17),
    .C1(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__o21a_1 _1741_ (.A1(net300),
    .A2(net14),
    .B1(_0471_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _1742_ (.A0(\lfsr0.seed_reg[20] ),
    .A1(\lfsr0.stop_reg[20] ),
    .S(net69),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _1743_ (.A1(_1267_),
    .A2(net41),
    .B1(_0472_),
    .B2(net62),
    .X(_0473_));
 sky130_fd_sc_hd__a211o_1 _1744_ (.A1(\sa0.signature_o[20] ),
    .A2(net20),
    .B1(net17),
    .C1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__o21a_1 _1745_ (.A1(net330),
    .A2(net14),
    .B1(_0474_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _1746_ (.A0(\lfsr0.seed_reg[21] ),
    .A1(\lfsr0.stop_reg[21] ),
    .S(net69),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _1747_ (.A1(_1239_),
    .A2(net40),
    .B1(_0475_),
    .B2(net60),
    .X(_0476_));
 sky130_fd_sc_hd__a211o_1 _1748_ (.A1(\sa0.signature_o[21] ),
    .A2(net20),
    .B1(net17),
    .C1(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__o21a_1 _1749_ (.A1(net313),
    .A2(net16),
    .B1(_0477_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _1750_ (.A0(\lfsr0.seed_reg[22] ),
    .A1(\lfsr0.stop_reg[22] ),
    .S(net69),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _1751_ (.A1(_1257_),
    .A2(net40),
    .B1(_0478_),
    .B2(net60),
    .X(_0479_));
 sky130_fd_sc_hd__a211o_1 _1752_ (.A1(\sa0.signature_o[22] ),
    .A2(net20),
    .B1(net17),
    .C1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__o21a_1 _1753_ (.A1(net301),
    .A2(net14),
    .B1(_0480_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _1754_ (.A0(\lfsr0.seed_reg[23] ),
    .A1(\lfsr0.stop_reg[23] ),
    .S(net69),
    .X(_0481_));
 sky130_fd_sc_hd__a22o_1 _1755_ (.A1(_1271_),
    .A2(net40),
    .B1(_0481_),
    .B2(net60),
    .X(_0482_));
 sky130_fd_sc_hd__a211o_1 _1756_ (.A1(\sa0.signature_o[23] ),
    .A2(net20),
    .B1(net17),
    .C1(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__o21a_1 _1757_ (.A1(net296),
    .A2(net14),
    .B1(_0483_),
    .X(_0173_));
 sky130_fd_sc_hd__a21oi_1 _1758_ (.A1(\sa0.en_i ),
    .A2(_0383_),
    .B1(\sa0.clear_i ),
    .Y(_0484_));
 sky130_fd_sc_hd__and3b_1 _1759_ (.A_N(\sa0.clear_i ),
    .B(_0383_),
    .C(\sa0.en_i ),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _1760_ (.A1(net456),
    .A2(net38),
    .B1(net35),
    .B2(_0391_),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _1761_ (.A(\sa0.signature_o[0] ),
    .B(_0397_),
    .Y(_0486_));
 sky130_fd_sc_hd__or2_1 _1762_ (.A(\sa0.signature_o[0] ),
    .B(_0397_),
    .X(_0487_));
 sky130_fd_sc_hd__a32o_1 _1763_ (.A1(net35),
    .A2(_0486_),
    .A3(_0487_),
    .B1(net38),
    .B2(net406),
    .X(_0175_));
 sky130_fd_sc_hd__nand2_1 _1764_ (.A(\sa0.signature_o[1] ),
    .B(_0403_),
    .Y(_0488_));
 sky130_fd_sc_hd__or2_1 _1765_ (.A(\sa0.signature_o[1] ),
    .B(_0403_),
    .X(_0489_));
 sky130_fd_sc_hd__a32o_1 _1766_ (.A1(net35),
    .A2(_0488_),
    .A3(_0489_),
    .B1(net38),
    .B2(net409),
    .X(_0176_));
 sky130_fd_sc_hd__nand2_1 _1767_ (.A(\sa0.signature_o[2] ),
    .B(_0409_),
    .Y(_0490_));
 sky130_fd_sc_hd__or2_1 _1768_ (.A(\sa0.signature_o[2] ),
    .B(_0409_),
    .X(_0491_));
 sky130_fd_sc_hd__a32o_1 _1769_ (.A1(net35),
    .A2(_0490_),
    .A3(_0491_),
    .B1(net38),
    .B2(net407),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _1770_ (.A(\sa0.signature_o[3] ),
    .B(_0414_),
    .Y(_0492_));
 sky130_fd_sc_hd__or2_1 _1771_ (.A(\sa0.signature_o[3] ),
    .B(_0414_),
    .X(_0493_));
 sky130_fd_sc_hd__a32o_1 _1772_ (.A1(net36),
    .A2(_0492_),
    .A3(_0493_),
    .B1(net39),
    .B2(net413),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _1773_ (.A(\sa0.signature_o[4] ),
    .B(_0419_),
    .Y(_0494_));
 sky130_fd_sc_hd__or2_1 _1774_ (.A(\sa0.signature_o[4] ),
    .B(_0419_),
    .X(_0495_));
 sky130_fd_sc_hd__a32o_1 _1775_ (.A1(net36),
    .A2(_0494_),
    .A3(_0495_),
    .B1(net39),
    .B2(net410),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _1776_ (.A(\sa0.signature_o[5] ),
    .B(_0424_),
    .Y(_0496_));
 sky130_fd_sc_hd__or2_1 _1777_ (.A(\sa0.signature_o[5] ),
    .B(_0424_),
    .X(_0497_));
 sky130_fd_sc_hd__a32o_1 _1778_ (.A1(net36),
    .A2(_0496_),
    .A3(_0497_),
    .B1(net39),
    .B2(net405),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _1779_ (.A(\sa0.signature_o[6] ),
    .B(_0429_),
    .Y(_0498_));
 sky130_fd_sc_hd__or2_1 _1780_ (.A(\sa0.signature_o[6] ),
    .B(_0429_),
    .X(_0499_));
 sky130_fd_sc_hd__a32o_1 _1781_ (.A1(net36),
    .A2(_0498_),
    .A3(_0499_),
    .B1(net39),
    .B2(net359),
    .X(_0181_));
 sky130_fd_sc_hd__a22o_1 _1782_ (.A1(net365),
    .A2(net39),
    .B1(net36),
    .B2(net359),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_1 _1783_ (.A1(net396),
    .A2(net37),
    .B1(net34),
    .B2(net365),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _1784_ (.A1(net385),
    .A2(net37),
    .B1(net34),
    .B2(net396),
    .X(_0184_));
 sky130_fd_sc_hd__a22o_1 _1785_ (.A1(net370),
    .A2(net37),
    .B1(net34),
    .B2(net385),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _1786_ (.A1(\sa0.signature_o[12] ),
    .A2(net38),
    .B1(net35),
    .B2(net370),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _1787_ (.A1(\sa0.signature_o[13] ),
    .A2(net37),
    .B1(net34),
    .B2(net400),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_1 _1788_ (.A1(net377),
    .A2(net37),
    .B1(net34),
    .B2(net404),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _1789_ (.A1(\sa0.signature_o[15] ),
    .A2(net37),
    .B1(net34),
    .B2(net377),
    .X(_0189_));
 sky130_fd_sc_hd__a22o_1 _1790_ (.A1(\sa0.signature_o[16] ),
    .A2(net38),
    .B1(net35),
    .B2(net380),
    .X(_0190_));
 sky130_fd_sc_hd__a22o_1 _1791_ (.A1(net360),
    .A2(net38),
    .B1(net35),
    .B2(net384),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _1792_ (.A1(\sa0.signature_o[18] ),
    .A2(net38),
    .B1(net35),
    .B2(net360),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_1 _1793_ (.A1(\sa0.signature_o[19] ),
    .A2(net38),
    .B1(net35),
    .B2(net382),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_1 _1794_ (.A1(\sa0.signature_o[20] ),
    .A2(net37),
    .B1(net34),
    .B2(net386),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _1795_ (.A1(net388),
    .A2(net37),
    .B1(net34),
    .B2(net392),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _1796_ (.A1(\sa0.signature_o[22] ),
    .A2(net37),
    .B1(net34),
    .B2(net388),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_1 _1797_ (.A1(net317),
    .A2(net37),
    .B1(net34),
    .B2(\sa0.signature_o[22] ),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _1798_ (.A(\gray_sobel0.sobel0.counter_sobel[1] ),
    .B(\gray_sobel0.sobel0.counter_sobel[0] ),
    .Y(_0500_));
 sky130_fd_sc_hd__o31a_1 _1799_ (.A1(\gray_sobel0.sobel0.counter_sobel[2] ),
    .A2(\gray_sobel0.sobel0.counter_sobel[3] ),
    .A3(_0500_),
    .B1(net33),
    .X(_0501_));
 sky130_fd_sc_hd__or4_4 _1800_ (.A(\gray_sobel0.sobel0.counter_sobel[2] ),
    .B(\gray_sobel0.sobel0.counter_sobel[3] ),
    .C(_1222_),
    .D(_1224_),
    .X(_0502_));
 sky130_fd_sc_hd__o21a_4 _1801_ (.A1(net47),
    .A2(_1222_),
    .B1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__nor2_4 _1802_ (.A(_0501_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__and2b_1 _1803_ (.A_N(net42),
    .B(_0390_),
    .X(_0505_));
 sky130_fd_sc_hd__a21o_1 _1804_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ),
    .A2(net42),
    .B1(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(net430),
    .A1(_0506_),
    .S(_0504_),
    .X(_0198_));
 sky130_fd_sc_hd__and2b_1 _1806_ (.A_N(net42),
    .B(_0396_),
    .X(_0507_));
 sky130_fd_sc_hd__a21o_1 _1807_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ),
    .A2(net43),
    .B1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1808_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[1] ),
    .A1(_0508_),
    .S(_0504_),
    .X(_0199_));
 sky130_fd_sc_hd__and2b_1 _1809_ (.A_N(net43),
    .B(_0402_),
    .X(_0509_));
 sky130_fd_sc_hd__a21o_1 _1810_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[2] ),
    .A2(net45),
    .B1(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _1811_ (.A0(net201),
    .A1(_0510_),
    .S(_0504_),
    .X(_0200_));
 sky130_fd_sc_hd__and2b_1 _1812_ (.A_N(net44),
    .B(_0408_),
    .X(_0511_));
 sky130_fd_sc_hd__a21o_1 _1813_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ),
    .A2(net44),
    .B1(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _1814_ (.A0(net416),
    .A1(_0512_),
    .S(_0504_),
    .X(_0201_));
 sky130_fd_sc_hd__and2b_1 _1815_ (.A_N(net45),
    .B(_0413_),
    .X(_0513_));
 sky130_fd_sc_hd__a21o_1 _1816_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ),
    .A2(net44),
    .B1(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _1817_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[4] ),
    .A1(_0514_),
    .S(_0504_),
    .X(_0202_));
 sky130_fd_sc_hd__and2b_2 _1818_ (.A_N(net46),
    .B(_0418_),
    .X(_0515_));
 sky130_fd_sc_hd__a21o_1 _1819_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ),
    .A2(net46),
    .B1(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _1820_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[5] ),
    .A1(_0516_),
    .S(_0504_),
    .X(_0203_));
 sky130_fd_sc_hd__and2b_1 _1821_ (.A_N(net49),
    .B(_0423_),
    .X(_0517_));
 sky130_fd_sc_hd__a21o_1 _1822_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[6] ),
    .A2(net49),
    .B1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _1823_ (.A0(net204),
    .A1(_0518_),
    .S(_0504_),
    .X(_0204_));
 sky130_fd_sc_hd__and2b_1 _1824_ (.A_N(net48),
    .B(_0428_),
    .X(_0519_));
 sky130_fd_sc_hd__a21o_1 _1825_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ),
    .A2(net48),
    .B1(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _1826_ (.A0(net403),
    .A1(_0520_),
    .S(_0504_),
    .X(_0205_));
 sky130_fd_sc_hd__nand2b_1 _1827_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[2] ),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2b_1 _1828_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[2] ),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _1829_ (.A(_0521_),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__and2b_1 _1830_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[1] ),
    .X(_0524_));
 sky130_fd_sc_hd__nand2b_1 _1831_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[0] ),
    .Y(_0525_));
 sky130_fd_sc_hd__xnor2_1 _1832_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[1] ),
    .Y(_0526_));
 sky130_fd_sc_hd__a21oi_1 _1833_ (.A1(_0525_),
    .A2(_0526_),
    .B1(_0524_),
    .Y(_0527_));
 sky130_fd_sc_hd__xnor2_1 _1834_ (.A(_0523_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2b_1 _1835_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2b_1 _1836_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[2] ),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1837_ (.A(_0529_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__and2b_1 _1838_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ),
    .X(_0532_));
 sky130_fd_sc_hd__nand2b_1 _1839_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ),
    .Y(_0533_));
 sky130_fd_sc_hd__xnor2_1 _1840_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ),
    .Y(_0534_));
 sky130_fd_sc_hd__a21oi_1 _1841_ (.A1(_0533_),
    .A2(_0534_),
    .B1(_0532_),
    .Y(_0535_));
 sky130_fd_sc_hd__o21ai_1 _1842_ (.A1(_0531_),
    .A2(_0535_),
    .B1(_0529_),
    .Y(_0536_));
 sky130_fd_sc_hd__and2b_1 _1843_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ),
    .X(_0537_));
 sky130_fd_sc_hd__nand2b_1 _1844_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ),
    .Y(_0538_));
 sky130_fd_sc_hd__and2b_1 _1845_ (.A_N(_0537_),
    .B(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__xnor2_1 _1846_ (.A(_0536_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nor2_1 _1847_ (.A(_0528_),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__xor2_1 _1848_ (.A(_0528_),
    .B(_0540_),
    .X(_0542_));
 sky130_fd_sc_hd__and2b_1 _1849_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[2] ),
    .X(_0543_));
 sky130_fd_sc_hd__and2b_1 _1850_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[2] ),
    .X(_0544_));
 sky130_fd_sc_hd__nor2_1 _1851_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__and2b_1 _1852_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[1] ),
    .X(_0546_));
 sky130_fd_sc_hd__nand2b_1 _1853_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[0] ),
    .Y(_0547_));
 sky130_fd_sc_hd__xnor2_2 _1854_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[1] ),
    .Y(_0548_));
 sky130_fd_sc_hd__a21oi_1 _1855_ (.A1(_0547_),
    .A2(_0548_),
    .B1(_0546_),
    .Y(_0549_));
 sky130_fd_sc_hd__o21bai_1 _1856_ (.A1(_0544_),
    .A2(_0549_),
    .B1_N(_0543_),
    .Y(_0550_));
 sky130_fd_sc_hd__nor2_1 _1857_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[3] ),
    .B(_1165_),
    .Y(_0551_));
 sky130_fd_sc_hd__and2_1 _1858_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[3] ),
    .B(_1165_),
    .X(_0552_));
 sky130_fd_sc_hd__nor2_1 _1859_ (.A(_0551_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__xor2_1 _1860_ (.A(_0550_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__xnor2_1 _1861_ (.A(_0542_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__xnor2_1 _1862_ (.A(_0525_),
    .B(_0526_),
    .Y(_0556_));
 sky130_fd_sc_hd__xnor2_1 _1863_ (.A(_0531_),
    .B(_0535_),
    .Y(_0557_));
 sky130_fd_sc_hd__nor2_1 _1864_ (.A(_0556_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__xnor2_1 _1865_ (.A(_0545_),
    .B(_0549_),
    .Y(_0559_));
 sky130_fd_sc_hd__xor2_1 _1866_ (.A(_0556_),
    .B(_0557_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _1867_ (.A1(_0559_),
    .A2(_0560_),
    .B1(_0558_),
    .Y(_0561_));
 sky130_fd_sc_hd__nor2_1 _1868_ (.A(_0555_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__xnor2_1 _1869_ (.A(_0559_),
    .B(_0560_),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2b_1 _1870_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[0] ),
    .Y(_0564_));
 sky130_fd_sc_hd__xnor2_1 _1871_ (.A(_0533_),
    .B(_0534_),
    .Y(_0565_));
 sky130_fd_sc_hd__a21oi_1 _1872_ (.A1(_0525_),
    .A2(_0564_),
    .B1(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__xor2_2 _1873_ (.A(_0547_),
    .B(_0548_),
    .X(_0567_));
 sky130_fd_sc_hd__and3_1 _1874_ (.A(_0525_),
    .B(_0564_),
    .C(_0565_),
    .X(_0568_));
 sky130_fd_sc_hd__nor2_1 _1875_ (.A(_0566_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__a21oi_1 _1876_ (.A1(_0567_),
    .A2(_0569_),
    .B1(_0566_),
    .Y(_0570_));
 sky130_fd_sc_hd__nor2_1 _1877_ (.A(_0563_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__xor2_1 _1878_ (.A(_0563_),
    .B(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__xor2_2 _1879_ (.A(_0567_),
    .B(_0569_),
    .X(_0573_));
 sky130_fd_sc_hd__nand2b_1 _1880_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ),
    .Y(_0574_));
 sky130_fd_sc_hd__xnor2_1 _1881_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[0] ),
    .Y(_0575_));
 sky130_fd_sc_hd__a21oi_1 _1882_ (.A1(_0533_),
    .A2(_0574_),
    .B1(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__and2_1 _1883_ (.A(_0573_),
    .B(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__a21o_1 _1884_ (.A1(_0572_),
    .A2(_0577_),
    .B1(_0571_),
    .X(_0578_));
 sky130_fd_sc_hd__xor2_1 _1885_ (.A(_0555_),
    .B(_0561_),
    .X(_0579_));
 sky130_fd_sc_hd__a21o_1 _1886_ (.A1(_0578_),
    .A2(_0579_),
    .B1(_0562_),
    .X(_0580_));
 sky130_fd_sc_hd__nand2b_1 _1887_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2b_1 _1888_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ),
    .Y(_0582_));
 sky130_fd_sc_hd__nand2_1 _1889_ (.A(_0581_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__a31oi_1 _1890_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ),
    .A2(_1161_),
    .A3(_0538_),
    .B1(_0537_),
    .Y(_0584_));
 sky130_fd_sc_hd__or3b_1 _1891_ (.A(_0531_),
    .B(_0535_),
    .C_N(_0539_),
    .X(_0585_));
 sky130_fd_sc_hd__a21o_1 _1892_ (.A1(_0584_),
    .A2(_0585_),
    .B1(_0583_),
    .X(_0586_));
 sky130_fd_sc_hd__nand3_1 _1893_ (.A(_0583_),
    .B(_0584_),
    .C(_0585_),
    .Y(_0587_));
 sky130_fd_sc_hd__o21ai_1 _1894_ (.A1(_0523_),
    .A2(_0527_),
    .B1(_0521_),
    .Y(_0588_));
 sky130_fd_sc_hd__and2b_1 _1895_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[3] ),
    .X(_0589_));
 sky130_fd_sc_hd__nand2b_1 _1896_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[3] ),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2b_1 _1897_ (.A_N(_0589_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__xnor2_1 _1898_ (.A(_0588_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__and3_1 _1899_ (.A(_0586_),
    .B(_0587_),
    .C(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__a21oi_1 _1900_ (.A1(_0586_),
    .A2(_0587_),
    .B1(_0592_),
    .Y(_0594_));
 sky130_fd_sc_hd__a21o_1 _1901_ (.A1(_0550_),
    .A2(_0553_),
    .B1(_0551_),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _1902_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[4] ),
    .B(_1164_),
    .Y(_0596_));
 sky130_fd_sc_hd__and2_1 _1903_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[4] ),
    .B(_1164_),
    .X(_0597_));
 sky130_fd_sc_hd__nor2_1 _1904_ (.A(_0596_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__xnor2_1 _1905_ (.A(_0595_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__or3_1 _1906_ (.A(_0593_),
    .B(_0594_),
    .C(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__o21ai_1 _1907_ (.A1(_0593_),
    .A2(_0594_),
    .B1(_0599_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2_1 _1908_ (.A(_0600_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__a21o_1 _1909_ (.A1(_0542_),
    .A2(_0554_),
    .B1(_0541_),
    .X(_0603_));
 sky130_fd_sc_hd__and3_1 _1910_ (.A(_0600_),
    .B(_0601_),
    .C(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__xnor2_1 _1911_ (.A(_0602_),
    .B(_0603_),
    .Y(_0605_));
 sky130_fd_sc_hd__xnor2_1 _1912_ (.A(_0580_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__xor2_1 _1913_ (.A(_0578_),
    .B(_0579_),
    .X(_0607_));
 sky130_fd_sc_hd__xnor2_1 _1914_ (.A(_0572_),
    .B(_0577_),
    .Y(_0608_));
 sky130_fd_sc_hd__and3_1 _1915_ (.A(_0533_),
    .B(_0574_),
    .C(_0575_),
    .X(_0609_));
 sky130_fd_sc_hd__nor2_2 _1916_ (.A(_0576_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__nor2_1 _1917_ (.A(_0573_),
    .B(_0576_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _1918_ (.A(_0577_),
    .B(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__nor2_1 _1919_ (.A(_0610_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__nand2_1 _1920_ (.A(_0608_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _1921_ (.A(_0607_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_1 _1922_ (.A(_0606_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a21o_1 _1923_ (.A1(_0588_),
    .A2(_0590_),
    .B1(_0589_),
    .X(_0617_));
 sky130_fd_sc_hd__and2b_1 _1924_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[4] ),
    .X(_0618_));
 sky130_fd_sc_hd__and2b_1 _1925_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[4] ),
    .X(_0619_));
 sky130_fd_sc_hd__nor2_1 _1926_ (.A(_0618_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__xnor2_1 _1927_ (.A(_0617_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__and2_1 _1928_ (.A(_1158_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_1 _1929_ (.A(_1158_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ),
    .Y(_0623_));
 sky130_fd_sc_hd__nor2_1 _1930_ (.A(_0622_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand3_1 _1931_ (.A(_0581_),
    .B(_0586_),
    .C(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__a21o_1 _1932_ (.A1(_0581_),
    .A2(_0586_),
    .B1(_0624_),
    .X(_0626_));
 sky130_fd_sc_hd__a21o_1 _1933_ (.A1(_0625_),
    .A2(_0626_),
    .B1(_0621_),
    .X(_0627_));
 sky130_fd_sc_hd__nand3_1 _1934_ (.A(_0621_),
    .B(_0625_),
    .C(_0626_),
    .Y(_0628_));
 sky130_fd_sc_hd__and2b_1 _1935_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[5] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[5] ),
    .X(_0629_));
 sky130_fd_sc_hd__nand2b_1 _1936_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[5] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[5] ),
    .Y(_0630_));
 sky130_fd_sc_hd__and2b_1 _1937_ (.A_N(_0629_),
    .B(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__a21oi_1 _1938_ (.A1(_0595_),
    .A2(_0598_),
    .B1(_0596_),
    .Y(_0632_));
 sky130_fd_sc_hd__xnor2_1 _1939_ (.A(_0631_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand3_1 _1940_ (.A(_0627_),
    .B(_0628_),
    .C(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__a21o_1 _1941_ (.A1(_0627_),
    .A2(_0628_),
    .B1(_0633_),
    .X(_0635_));
 sky130_fd_sc_hd__nand2b_1 _1942_ (.A_N(_0593_),
    .B(_0600_),
    .Y(_0636_));
 sky130_fd_sc_hd__a21oi_1 _1943_ (.A1(_0634_),
    .A2(_0635_),
    .B1(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21o_1 _1944_ (.A1(_0634_),
    .A2(_0635_),
    .B1(_0636_),
    .X(_0638_));
 sky130_fd_sc_hd__and3_1 _1945_ (.A(_0634_),
    .B(_0635_),
    .C(_0636_),
    .X(_0639_));
 sky130_fd_sc_hd__or2_1 _1946_ (.A(_0637_),
    .B(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__a21o_1 _1947_ (.A1(_0580_),
    .A2(_0605_),
    .B1(_0604_),
    .X(_0641_));
 sky130_fd_sc_hd__xnor2_1 _1948_ (.A(_0640_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nor2_1 _1949_ (.A(_0616_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__xor2_1 _1950_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[6] ),
    .X(_0644_));
 sky130_fd_sc_hd__inv_2 _1951_ (.A(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21a_1 _1952_ (.A1(_1158_),
    .A2(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ),
    .B1(_0581_),
    .X(_0646_));
 sky130_fd_sc_hd__a21oi_1 _1953_ (.A1(_0586_),
    .A2(_0646_),
    .B1(_0622_),
    .Y(_0647_));
 sky130_fd_sc_hd__xnor2_1 _1954_ (.A(_0644_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__xnor2_1 _1955_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[5] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[5] ),
    .Y(_0649_));
 sky130_fd_sc_hd__a21oi_1 _1956_ (.A1(_0617_),
    .A2(_0620_),
    .B1(_0618_),
    .Y(_0650_));
 sky130_fd_sc_hd__xnor2_1 _1957_ (.A(_0649_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__and2_1 _1958_ (.A(_0648_),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__xor2_1 _1959_ (.A(_0648_),
    .B(_0651_),
    .X(_0653_));
 sky130_fd_sc_hd__and2b_1 _1960_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[6] ),
    .X(_0654_));
 sky130_fd_sc_hd__nand2b_1 _1961_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[6] ),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2b_1 _1962_ (.A_N(_0654_),
    .B(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21oi_1 _1963_ (.A1(_0630_),
    .A2(_0632_),
    .B1(_0629_),
    .Y(_0657_));
 sky130_fd_sc_hd__xnor2_1 _1964_ (.A(_0656_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__xnor2_1 _1965_ (.A(_0653_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__and2_1 _1966_ (.A(_0627_),
    .B(_0634_),
    .X(_0660_));
 sky130_fd_sc_hd__nor2_1 _1967_ (.A(_0659_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__xor2_1 _1968_ (.A(_0659_),
    .B(_0660_),
    .X(_0662_));
 sky130_fd_sc_hd__a211o_1 _1969_ (.A1(_0580_),
    .A2(_0605_),
    .B1(_0639_),
    .C1(_0604_),
    .X(_0663_));
 sky130_fd_sc_hd__and3_1 _1970_ (.A(_0638_),
    .B(_0662_),
    .C(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__a21oi_1 _1971_ (.A1(_0638_),
    .A2(_0663_),
    .B1(_0662_),
    .Y(_0665_));
 sky130_fd_sc_hd__or2_1 _1972_ (.A(_0664_),
    .B(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__nand2_1 _1973_ (.A(_0643_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__and2b_1 _1974_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[7] ),
    .X(_0668_));
 sky130_fd_sc_hd__nand2b_1 _1975_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[7] ),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2b_1 _1976_ (.A_N(_0668_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__a21o_1 _1977_ (.A1(_0655_),
    .A2(_0657_),
    .B1(_0654_),
    .X(_0671_));
 sky130_fd_sc_hd__a21oi_2 _1978_ (.A1(_0669_),
    .A2(_0671_),
    .B1(_0668_),
    .Y(_0672_));
 sky130_fd_sc_hd__and2b_1 _1979_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ),
    .X(_0673_));
 sky130_fd_sc_hd__a22o_1 _1980_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ),
    .A2(_1162_),
    .B1(_0645_),
    .B2(_0647_),
    .X(_0674_));
 sky130_fd_sc_hd__and2b_1 _1981_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _1982_ (.A(_0673_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__a21oi_2 _1983_ (.A1(_0674_),
    .A2(_0676_),
    .B1(_0673_),
    .Y(_0677_));
 sky130_fd_sc_hd__and2b_1 _1984_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[7] ),
    .X(_0678_));
 sky130_fd_sc_hd__nand2b_1 _1985_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[7] ),
    .Y(_0679_));
 sky130_fd_sc_hd__nand2b_1 _1986_ (.A_N(_0678_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__and2b_1 _1987_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[6] ),
    .X(_0681_));
 sky130_fd_sc_hd__nand2b_1 _1988_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[6] ),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2b_1 _1989_ (.A_N(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a21oi_1 _1990_ (.A1(_1163_),
    .A2(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[5] ),
    .B1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[4] ),
    .Y(_0684_));
 sky130_fd_sc_hd__a2bb2o_1 _1991_ (.A1_N(_1163_),
    .A2_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[5] ),
    .B1(_0684_),
    .B2(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[4] ),
    .X(_0685_));
 sky130_fd_sc_hd__a31o_1 _1992_ (.A1(_0617_),
    .A2(_0620_),
    .A3(_0649_),
    .B1(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__a21o_1 _1993_ (.A1(_0682_),
    .A2(_0686_),
    .B1(_0681_),
    .X(_0687_));
 sky130_fd_sc_hd__a21oi_1 _1994_ (.A1(_0679_),
    .A2(_0687_),
    .B1(_0678_),
    .Y(_0688_));
 sky130_fd_sc_hd__nor2_1 _1995_ (.A(_0677_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__or3_4 _1996_ (.A(_0672_),
    .B(_0677_),
    .C(_0688_),
    .X(_0690_));
 sky130_fd_sc_hd__xnor2_1 _1997_ (.A(_0680_),
    .B(_0687_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand2_1 _1998_ (.A(_0677_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__xor2_1 _1999_ (.A(_0677_),
    .B(_0691_),
    .X(_0693_));
 sky130_fd_sc_hd__nand2_1 _2000_ (.A(_0672_),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__and2_1 _2001_ (.A(_0677_),
    .B(_0688_),
    .X(_0695_));
 sky130_fd_sc_hd__nor2_1 _2002_ (.A(_0689_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__xnor2_1 _2003_ (.A(_0672_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a21oi_1 _2004_ (.A1(_0692_),
    .A2(_0694_),
    .B1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a21o_1 _2005_ (.A1(_0692_),
    .A2(_0694_),
    .B1(_0697_),
    .X(_0699_));
 sky130_fd_sc_hd__or2_1 _2006_ (.A(_0672_),
    .B(_0693_),
    .X(_0700_));
 sky130_fd_sc_hd__nand2_1 _2007_ (.A(_0694_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__xor2_1 _2008_ (.A(_0674_),
    .B(_0676_),
    .X(_0702_));
 sky130_fd_sc_hd__xnor2_1 _2009_ (.A(_0683_),
    .B(_0686_),
    .Y(_0703_));
 sky130_fd_sc_hd__and2_1 _2010_ (.A(_0702_),
    .B(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__xor2_1 _2011_ (.A(_0702_),
    .B(_0703_),
    .X(_0705_));
 sky130_fd_sc_hd__xnor2_1 _2012_ (.A(_0670_),
    .B(_0671_),
    .Y(_0706_));
 sky130_fd_sc_hd__a21oi_1 _2013_ (.A1(_0705_),
    .A2(_0706_),
    .B1(_0704_),
    .Y(_0707_));
 sky130_fd_sc_hd__or2_1 _2014_ (.A(_0701_),
    .B(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__xnor2_1 _2015_ (.A(_0705_),
    .B(_0706_),
    .Y(_0709_));
 sky130_fd_sc_hd__a21oi_1 _2016_ (.A1(_0653_),
    .A2(_0658_),
    .B1(_0652_),
    .Y(_0710_));
 sky130_fd_sc_hd__nor2_1 _2017_ (.A(_0709_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__xor2_1 _2018_ (.A(_0709_),
    .B(_0710_),
    .X(_0712_));
 sky130_fd_sc_hd__a31o_1 _2019_ (.A1(_0638_),
    .A2(_0662_),
    .A3(_0663_),
    .B1(_0661_),
    .X(_0713_));
 sky130_fd_sc_hd__a21oi_1 _2020_ (.A1(_0712_),
    .A2(_0713_),
    .B1(_0711_),
    .Y(_0714_));
 sky130_fd_sc_hd__xnor2_1 _2021_ (.A(_0701_),
    .B(_0707_),
    .Y(_0715_));
 sky130_fd_sc_hd__o21a_1 _2022_ (.A1(_0714_),
    .A2(_0715_),
    .B1(_0708_),
    .X(_0716_));
 sky130_fd_sc_hd__o211a_2 _2023_ (.A1(_0714_),
    .A2(_0715_),
    .B1(_0699_),
    .C1(_0708_),
    .X(_0717_));
 sky130_fd_sc_hd__and3_1 _2024_ (.A(_0692_),
    .B(_0694_),
    .C(_0697_),
    .X(_0718_));
 sky130_fd_sc_hd__a21o_2 _2025_ (.A1(_0672_),
    .A2(_0695_),
    .B1(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__o21a_1 _2026_ (.A1(_0717_),
    .A2(_0719_),
    .B1(_0690_),
    .X(_0720_));
 sky130_fd_sc_hd__o21ai_2 _2027_ (.A1(_0717_),
    .A2(_0719_),
    .B1(_0690_),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_1 _2028_ (.A(_0667_),
    .B(_0720_),
    .Y(_0722_));
 sky130_fd_sc_hd__xor2_1 _2029_ (.A(_0712_),
    .B(_0713_),
    .X(_0723_));
 sky130_fd_sc_hd__xor2_1 _2030_ (.A(_0722_),
    .B(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__nand2b_1 _2031_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[2] ),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2b_1 _2032_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[2] ),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_1 _2033_ (.A(_0725_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__and2b_1 _2034_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[1] ),
    .X(_0728_));
 sky130_fd_sc_hd__nand2b_2 _2035_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[0] ),
    .Y(_0729_));
 sky130_fd_sc_hd__xnor2_1 _2036_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[1] ),
    .Y(_0730_));
 sky130_fd_sc_hd__a21oi_1 _2037_ (.A1(_0729_),
    .A2(_0730_),
    .B1(_0728_),
    .Y(_0731_));
 sky130_fd_sc_hd__xnor2_1 _2038_ (.A(_0727_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__or2_2 _2039_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ),
    .B(_1165_),
    .X(_0733_));
 sky130_fd_sc_hd__nand2_1 _2040_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ),
    .B(_1165_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _2041_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__and2b_1 _2042_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ),
    .X(_0736_));
 sky130_fd_sc_hd__nand2b_1 _2043_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[2] ),
    .Y(_0737_));
 sky130_fd_sc_hd__and2b_1 _2044_ (.A_N(_0736_),
    .B(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__and2b_1 _2045_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ),
    .X(_0739_));
 sky130_fd_sc_hd__nand2b_1 _2046_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[0] ),
    .Y(_0740_));
 sky130_fd_sc_hd__xnor2_1 _2047_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[1] ),
    .Y(_0741_));
 sky130_fd_sc_hd__a21o_1 _2048_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0739_),
    .X(_0742_));
 sky130_fd_sc_hd__a21oi_1 _2049_ (.A1(_0737_),
    .A2(_0742_),
    .B1(_0736_),
    .Y(_0743_));
 sky130_fd_sc_hd__xnor2_1 _2050_ (.A(_0735_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__nor2_1 _2051_ (.A(_0732_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__xor2_1 _2052_ (.A(_0732_),
    .B(_0744_),
    .X(_0746_));
 sky130_fd_sc_hd__nor2_1 _2053_ (.A(_1161_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[2] ),
    .Y(_0747_));
 sky130_fd_sc_hd__and2_1 _2054_ (.A(_1161_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[2] ),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_1 _2055_ (.A(_0747_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__and2b_1 _2056_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ),
    .X(_0750_));
 sky130_fd_sc_hd__nand2b_1 _2057_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[0] ),
    .Y(_0751_));
 sky130_fd_sc_hd__xnor2_1 _2058_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[1] ),
    .Y(_0752_));
 sky130_fd_sc_hd__a21oi_1 _2059_ (.A1(_0751_),
    .A2(_0752_),
    .B1(_0750_),
    .Y(_0753_));
 sky130_fd_sc_hd__o21bai_1 _2060_ (.A1(_0748_),
    .A2(_0753_),
    .B1_N(_0747_),
    .Y(_0754_));
 sky130_fd_sc_hd__and2b_1 _2061_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ),
    .X(_0755_));
 sky130_fd_sc_hd__and2b_1 _2062_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[3] ),
    .X(_0756_));
 sky130_fd_sc_hd__nor2_1 _2063_ (.A(_0755_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__xor2_1 _2064_ (.A(_0754_),
    .B(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__xnor2_1 _2065_ (.A(_0746_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__xor2_1 _2066_ (.A(_0729_),
    .B(_0730_),
    .X(_0760_));
 sky130_fd_sc_hd__xor2_1 _2067_ (.A(_0738_),
    .B(_0742_),
    .X(_0761_));
 sky130_fd_sc_hd__and2_1 _2068_ (.A(_0760_),
    .B(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__xnor2_1 _2069_ (.A(_0749_),
    .B(_0753_),
    .Y(_0763_));
 sky130_fd_sc_hd__xor2_1 _2070_ (.A(_0760_),
    .B(_0761_),
    .X(_0764_));
 sky130_fd_sc_hd__a21oi_1 _2071_ (.A1(_0763_),
    .A2(_0764_),
    .B1(_0762_),
    .Y(_0765_));
 sky130_fd_sc_hd__nor2_1 _2072_ (.A(_0759_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__xnor2_1 _2073_ (.A(_0763_),
    .B(_0764_),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2b_1 _2074_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[0] ),
    .Y(_0768_));
 sky130_fd_sc_hd__xnor2_1 _2075_ (.A(_0740_),
    .B(_0741_),
    .Y(_0769_));
 sky130_fd_sc_hd__a21oi_1 _2076_ (.A1(_0729_),
    .A2(_0768_),
    .B1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__xor2_1 _2077_ (.A(_0751_),
    .B(_0752_),
    .X(_0771_));
 sky130_fd_sc_hd__and3_1 _2078_ (.A(_0729_),
    .B(_0768_),
    .C(_0769_),
    .X(_0772_));
 sky130_fd_sc_hd__nor2_1 _2079_ (.A(_0770_),
    .B(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__a21oi_1 _2080_ (.A1(_0771_),
    .A2(_0773_),
    .B1(_0770_),
    .Y(_0774_));
 sky130_fd_sc_hd__nor2_1 _2081_ (.A(_0767_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__xor2_1 _2082_ (.A(_0767_),
    .B(_0774_),
    .X(_0776_));
 sky130_fd_sc_hd__nand2b_1 _2083_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ),
    .Y(_0777_));
 sky130_fd_sc_hd__nand2b_1 _2084_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[0] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ),
    .Y(_0778_));
 sky130_fd_sc_hd__a22o_1 _2085_ (.A1(_0740_),
    .A2(_0777_),
    .B1(_0778_),
    .B2(_0751_),
    .X(_0779_));
 sky130_fd_sc_hd__xor2_1 _2086_ (.A(_0771_),
    .B(_0773_),
    .X(_0780_));
 sky130_fd_sc_hd__and2b_1 _2087_ (.A_N(_0779_),
    .B(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__a21o_1 _2088_ (.A1(_0776_),
    .A2(_0781_),
    .B1(_0775_),
    .X(_0782_));
 sky130_fd_sc_hd__xor2_1 _2089_ (.A(_0759_),
    .B(_0765_),
    .X(_0783_));
 sky130_fd_sc_hd__a21o_1 _2090_ (.A1(_0782_),
    .A2(_0783_),
    .B1(_0766_),
    .X(_0784_));
 sky130_fd_sc_hd__xnor2_2 _2091_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[4] ),
    .Y(_0785_));
 sky130_fd_sc_hd__a221o_2 _2092_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ),
    .A2(_1165_),
    .B1(_0737_),
    .B2(_0742_),
    .C1(_0736_),
    .X(_0786_));
 sky130_fd_sc_hd__nand2_1 _2093_ (.A(_0733_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__xnor2_1 _2094_ (.A(_0785_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__o21ai_1 _2095_ (.A1(_0727_),
    .A2(_0731_),
    .B1(_0725_),
    .Y(_0789_));
 sky130_fd_sc_hd__and2b_1 _2096_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[3] ),
    .X(_0790_));
 sky130_fd_sc_hd__and2b_1 _2097_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[3] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[3] ),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_1 _2098_ (.A(_0790_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__xor2_1 _2099_ (.A(_0789_),
    .B(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _2100_ (.A(_0788_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__xor2_1 _2101_ (.A(_0788_),
    .B(_0793_),
    .X(_0795_));
 sky130_fd_sc_hd__a21o_1 _2102_ (.A1(_0754_),
    .A2(_0757_),
    .B1(_0755_),
    .X(_0796_));
 sky130_fd_sc_hd__and2b_1 _2103_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ),
    .X(_0797_));
 sky130_fd_sc_hd__and2b_1 _2104_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[4] ),
    .X(_0798_));
 sky130_fd_sc_hd__nor2_1 _2105_ (.A(_0797_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__xor2_1 _2106_ (.A(_0796_),
    .B(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__nand2_1 _2107_ (.A(_0795_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__xnor2_1 _2108_ (.A(_0795_),
    .B(_0800_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21oi_1 _2109_ (.A1(_0746_),
    .A2(_0758_),
    .B1(_0745_),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_1 _2110_ (.A(_0802_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__xor2_1 _2111_ (.A(_0802_),
    .B(_0803_),
    .X(_0805_));
 sky130_fd_sc_hd__xnor2_1 _2112_ (.A(_0784_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__xor2_1 _2113_ (.A(_0782_),
    .B(_0783_),
    .X(_0807_));
 sky130_fd_sc_hd__xnor2_1 _2114_ (.A(_0776_),
    .B(_0781_),
    .Y(_0808_));
 sky130_fd_sc_hd__xor2_1 _2115_ (.A(_0779_),
    .B(_0780_),
    .X(_0809_));
 sky130_fd_sc_hd__and2b_1 _2116_ (.A_N(_0610_),
    .B(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_1 _2117_ (.A(_0808_),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__nor2_1 _2118_ (.A(_0807_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__nand2_1 _2119_ (.A(_0806_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a21o_1 _2120_ (.A1(_0789_),
    .A2(_0792_),
    .B1(_0790_),
    .X(_0814_));
 sky130_fd_sc_hd__and2b_1 _2121_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[4] ),
    .X(_0815_));
 sky130_fd_sc_hd__and2b_1 _2122_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[4] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[4] ),
    .X(_0816_));
 sky130_fd_sc_hd__nor2_1 _2123_ (.A(_0815_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__xor2_1 _2124_ (.A(_0814_),
    .B(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__and2_1 _2125_ (.A(_1158_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[5] ),
    .X(_0819_));
 sky130_fd_sc_hd__or2_1 _2126_ (.A(_1158_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[5] ),
    .X(_0820_));
 sky130_fd_sc_hd__nand2b_1 _2127_ (.A_N(_0819_),
    .B(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__a32o_1 _2128_ (.A1(_0733_),
    .A2(_0785_),
    .A3(_0786_),
    .B1(_1164_),
    .B2(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ),
    .X(_0822_));
 sky130_fd_sc_hd__xnor2_1 _2129_ (.A(_0821_),
    .B(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__and2_1 _2130_ (.A(_0818_),
    .B(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__nor2_1 _2131_ (.A(_0818_),
    .B(_0823_),
    .Y(_0825_));
 sky130_fd_sc_hd__nor2_1 _2132_ (.A(_0824_),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__and2b_1 _2133_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[5] ),
    .X(_0827_));
 sky130_fd_sc_hd__inv_2 _2134_ (.A(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__and2b_1 _2135_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[5] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ),
    .X(_0829_));
 sky130_fd_sc_hd__nor2_1 _2136_ (.A(_0827_),
    .B(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__a21oi_1 _2137_ (.A1(_0796_),
    .A2(_0799_),
    .B1(_0797_),
    .Y(_0831_));
 sky130_fd_sc_hd__xnor2_1 _2138_ (.A(_0830_),
    .B(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__xnor2_1 _2139_ (.A(_0826_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__and3_1 _2140_ (.A(_0794_),
    .B(_0801_),
    .C(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__a21o_1 _2141_ (.A1(_0794_),
    .A2(_0801_),
    .B1(_0833_),
    .X(_0835_));
 sky130_fd_sc_hd__and2b_1 _2142_ (.A_N(_0834_),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__a21oi_2 _2143_ (.A1(_0784_),
    .A2(_0805_),
    .B1(_0804_),
    .Y(_0837_));
 sky130_fd_sc_hd__xnor2_1 _2144_ (.A(_0836_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_1 _2145_ (.A(_0813_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__xor2_2 _2146_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[6] ),
    .X(_0840_));
 sky130_fd_sc_hd__a21bo_1 _2147_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ),
    .A2(_1164_),
    .B1_N(_0820_),
    .X(_0841_));
 sky130_fd_sc_hd__a31oi_4 _2148_ (.A1(_0733_),
    .A2(_0785_),
    .A3(_0786_),
    .B1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__nor2_1 _2149_ (.A(_0819_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__xor2_1 _2150_ (.A(_0840_),
    .B(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__xnor2_1 _2151_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[5] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[5] ),
    .Y(_0845_));
 sky130_fd_sc_hd__a21oi_1 _2152_ (.A1(_0814_),
    .A2(_0817_),
    .B1(_0815_),
    .Y(_0846_));
 sky130_fd_sc_hd__xnor2_1 _2153_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__and2b_1 _2154_ (.A_N(_0844_),
    .B(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__xnor2_1 _2155_ (.A(_0844_),
    .B(_0847_),
    .Y(_0849_));
 sky130_fd_sc_hd__nor2_1 _2156_ (.A(_1162_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[6] ),
    .Y(_0850_));
 sky130_fd_sc_hd__and2_1 _2157_ (.A(_1162_),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[6] ),
    .X(_0851_));
 sky130_fd_sc_hd__inv_2 _2158_ (.A(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__nor2_1 _2159_ (.A(_0850_),
    .B(_0851_),
    .Y(_0853_));
 sky130_fd_sc_hd__a211o_1 _2160_ (.A1(_0796_),
    .A2(_0799_),
    .B1(_0829_),
    .C1(_0797_),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _2161_ (.A(_0828_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__xnor2_1 _2162_ (.A(_0853_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__xnor2_1 _2163_ (.A(_0849_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__a21oi_1 _2164_ (.A1(_0826_),
    .A2(_0832_),
    .B1(_0824_),
    .Y(_0858_));
 sky130_fd_sc_hd__xnor2_1 _2165_ (.A(_0857_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__a21o_1 _2166_ (.A1(_0835_),
    .A2(_0837_),
    .B1(_0834_),
    .X(_0860_));
 sky130_fd_sc_hd__or2_1 _2167_ (.A(_0859_),
    .B(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__nand2_1 _2168_ (.A(_0859_),
    .B(_0860_),
    .Y(_0862_));
 sky130_fd_sc_hd__nand2_1 _2169_ (.A(_0861_),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__and2_1 _2170_ (.A(_0839_),
    .B(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__nand2b_1 _2171_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ),
    .Y(_0865_));
 sky130_fd_sc_hd__xnor2_1 _2172_ (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[7] ),
    .Y(_0866_));
 sky130_fd_sc_hd__a31o_1 _2173_ (.A1(_0828_),
    .A2(_0852_),
    .A3(_0854_),
    .B1(_0850_),
    .X(_0867_));
 sky130_fd_sc_hd__nand2_1 _2174_ (.A(_0866_),
    .B(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand2_2 _2175_ (.A(_0865_),
    .B(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__and2b_1 _2176_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ),
    .X(_0870_));
 sky130_fd_sc_hd__o32ai_4 _2177_ (.A1(_0819_),
    .A2(_0840_),
    .A3(_0842_),
    .B1(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[6] ),
    .B2(_1159_),
    .Y(_0871_));
 sky130_fd_sc_hd__and2b_1 _2178_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[7] ),
    .X(_0872_));
 sky130_fd_sc_hd__nor2_1 _2179_ (.A(_0870_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21oi_2 _2180_ (.A1(_0871_),
    .A2(_0873_),
    .B1(_0870_),
    .Y(_0874_));
 sky130_fd_sc_hd__nand2b_1 _2181_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[7] ),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2b_1 _2182_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[7] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[7] ),
    .Y(_0876_));
 sky130_fd_sc_hd__nand2_1 _2183_ (.A(_0875_),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__and2b_1 _2184_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[6] ),
    .X(_0878_));
 sky130_fd_sc_hd__and2b_1 _2185_ (.A_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[6] ),
    .B(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[6] ),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_1 _2186_ (.A(_0878_),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__a21oi_1 _2187_ (.A1(_1160_),
    .A2(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[5] ),
    .B1(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[4] ),
    .Y(_0881_));
 sky130_fd_sc_hd__a2bb2o_1 _2188_ (.A1_N(_1160_),
    .A2_N(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[5] ),
    .B1(_0881_),
    .B2(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[4] ),
    .X(_0882_));
 sky130_fd_sc_hd__a31o_1 _2189_ (.A1(_0814_),
    .A2(_0817_),
    .A3(_0845_),
    .B1(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__a21oi_1 _2190_ (.A1(_0880_),
    .A2(_0883_),
    .B1(_0878_),
    .Y(_0884_));
 sky130_fd_sc_hd__or2_1 _2191_ (.A(_0877_),
    .B(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__and3_1 _2192_ (.A(_0874_),
    .B(_0875_),
    .C(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__xor2_1 _2193_ (.A(_0877_),
    .B(_0884_),
    .X(_0887_));
 sky130_fd_sc_hd__nand2_1 _2194_ (.A(_0874_),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__xor2_1 _2195_ (.A(_0874_),
    .B(_0887_),
    .X(_0889_));
 sky130_fd_sc_hd__nand2b_1 _2196_ (.A_N(_0869_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__a21oi_1 _2197_ (.A1(_0875_),
    .A2(_0885_),
    .B1(_0874_),
    .Y(_0891_));
 sky130_fd_sc_hd__or2_1 _2198_ (.A(_0886_),
    .B(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__xnor2_1 _2199_ (.A(_0869_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__and3_1 _2200_ (.A(_0888_),
    .B(_0890_),
    .C(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__xor2_1 _2201_ (.A(_0869_),
    .B(_0889_),
    .X(_0895_));
 sky130_fd_sc_hd__xnor2_1 _2202_ (.A(_0871_),
    .B(_0873_),
    .Y(_0896_));
 sky130_fd_sc_hd__xnor2_1 _2203_ (.A(_0880_),
    .B(_0883_),
    .Y(_0897_));
 sky130_fd_sc_hd__nor2_1 _2204_ (.A(_0896_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__xor2_1 _2205_ (.A(_0896_),
    .B(_0897_),
    .X(_0899_));
 sky130_fd_sc_hd__xor2_1 _2206_ (.A(_0866_),
    .B(_0867_),
    .X(_0900_));
 sky130_fd_sc_hd__a21oi_1 _2207_ (.A1(_0899_),
    .A2(_0900_),
    .B1(_0898_),
    .Y(_0901_));
 sky130_fd_sc_hd__or2_1 _2208_ (.A(_0895_),
    .B(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__xnor2_1 _2209_ (.A(_0899_),
    .B(_0900_),
    .Y(_0903_));
 sky130_fd_sc_hd__a21oi_1 _2210_ (.A1(_0849_),
    .A2(_0856_),
    .B1(_0848_),
    .Y(_0904_));
 sky130_fd_sc_hd__or2_1 _2211_ (.A(_0903_),
    .B(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__xnor2_1 _2212_ (.A(_0903_),
    .B(_0904_),
    .Y(_0906_));
 sky130_fd_sc_hd__a2111o_1 _2213_ (.A1(_0835_),
    .A2(_0837_),
    .B1(_0859_),
    .C1(_0906_),
    .D1(_0834_),
    .X(_0907_));
 sky130_fd_sc_hd__o31a_1 _2214_ (.A1(_0857_),
    .A2(_0858_),
    .A3(_0906_),
    .B1(_0905_),
    .X(_0908_));
 sky130_fd_sc_hd__xnor2_1 _2215_ (.A(_0895_),
    .B(_0901_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21o_1 _2216_ (.A1(_0907_),
    .A2(_0908_),
    .B1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__nand2_1 _2217_ (.A(_0902_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__and2_1 _2218_ (.A(_0869_),
    .B(_0891_),
    .X(_0912_));
 sky130_fd_sc_hd__nand2_2 _2219_ (.A(_0869_),
    .B(_0891_),
    .Y(_0913_));
 sky130_fd_sc_hd__a21o_1 _2220_ (.A1(_0888_),
    .A2(_0890_),
    .B1(_0893_),
    .X(_0914_));
 sky130_fd_sc_hd__a31o_1 _2221_ (.A1(_0865_),
    .A2(_0868_),
    .A3(_0886_),
    .B1(_0912_),
    .X(_0915_));
 sky130_fd_sc_hd__a311o_2 _2222_ (.A1(_0902_),
    .A2(_0910_),
    .A3(_0914_),
    .B1(_0915_),
    .C1(_0894_),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _2223_ (.A(_0913_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__or2_1 _2224_ (.A(_0864_),
    .B(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__o21a_1 _2225_ (.A1(_0857_),
    .A2(_0858_),
    .B1(_0861_),
    .X(_0919_));
 sky130_fd_sc_hd__xnor2_1 _2226_ (.A(_0906_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__xnor2_1 _2227_ (.A(_0918_),
    .B(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__nand2_1 _2228_ (.A(_0724_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__xor2_1 _2229_ (.A(_0714_),
    .B(_0715_),
    .X(_0923_));
 sky130_fd_sc_hd__nor2_1 _2230_ (.A(_0698_),
    .B(_0718_),
    .Y(_0924_));
 sky130_fd_sc_hd__xnor2_1 _2231_ (.A(_0716_),
    .B(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__o21a_1 _2232_ (.A1(_0923_),
    .A2(_0925_),
    .B1(_0721_),
    .X(_0926_));
 sky130_fd_sc_hd__and2b_1 _2233_ (.A_N(_0894_),
    .B(_0914_),
    .X(_0927_));
 sky130_fd_sc_hd__xnor2_1 _2234_ (.A(_0911_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand3_1 _2235_ (.A(_0907_),
    .B(_0908_),
    .C(_0909_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand2_1 _2236_ (.A(_0910_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand3_1 _2237_ (.A(_0917_),
    .B(_0928_),
    .C(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__a2111o_1 _2238_ (.A1(_0864_),
    .A2(_0920_),
    .B1(_0928_),
    .C1(_0930_),
    .D1(_0917_),
    .X(_0932_));
 sky130_fd_sc_hd__o211ai_1 _2239_ (.A1(_0667_),
    .A2(_0723_),
    .B1(_0923_),
    .C1(_0925_),
    .Y(_0933_));
 sky130_fd_sc_hd__a221o_1 _2240_ (.A1(_0931_),
    .A2(_0932_),
    .B1(_0933_),
    .B2(_0720_),
    .C1(_0926_),
    .X(_0934_));
 sky130_fd_sc_hd__and2_1 _2241_ (.A(_0616_),
    .B(_0720_),
    .X(_0935_));
 sky130_fd_sc_hd__xnor2_1 _2242_ (.A(_0642_),
    .B(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__and3_1 _2243_ (.A(_0813_),
    .B(_0913_),
    .C(_0916_),
    .X(_0937_));
 sky130_fd_sc_hd__xnor2_1 _2244_ (.A(_0838_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__nor2_1 _2245_ (.A(_0936_),
    .B(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__nor2_1 _2246_ (.A(_0615_),
    .B(_0721_),
    .Y(_0940_));
 sky130_fd_sc_hd__xor2_1 _2247_ (.A(_0606_),
    .B(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__or2_1 _2248_ (.A(_0812_),
    .B(_0917_),
    .X(_0942_));
 sky130_fd_sc_hd__xnor2_1 _2249_ (.A(_0806_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__nor2_1 _2250_ (.A(_0941_),
    .B(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__nand2_1 _2251_ (.A(_0941_),
    .B(_0943_),
    .Y(_0945_));
 sky130_fd_sc_hd__nand2b_1 _2252_ (.A_N(_0944_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__o211a_1 _2253_ (.A1(_0717_),
    .A2(_0719_),
    .B1(_0614_),
    .C1(_0690_),
    .X(_0947_));
 sky130_fd_sc_hd__xor2_1 _2254_ (.A(_0607_),
    .B(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__and3_1 _2255_ (.A(_0811_),
    .B(_0913_),
    .C(_0916_),
    .X(_0949_));
 sky130_fd_sc_hd__xor2_1 _2256_ (.A(_0807_),
    .B(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__nor2_1 _2257_ (.A(_0948_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__or2_1 _2258_ (.A(_0948_),
    .B(_0950_),
    .X(_0952_));
 sky130_fd_sc_hd__and2_1 _2259_ (.A(_0948_),
    .B(_0950_),
    .X(_0953_));
 sky130_fd_sc_hd__o221a_1 _2260_ (.A1(_0610_),
    .A2(_0612_),
    .B1(_0717_),
    .B2(_0719_),
    .C1(_0690_),
    .X(_0954_));
 sky130_fd_sc_hd__xnor2_1 _2261_ (.A(_0608_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__or3b_1 _2262_ (.A(_0810_),
    .B(_0912_),
    .C_N(_0916_),
    .X(_0956_));
 sky130_fd_sc_hd__xor2_1 _2263_ (.A(_0808_),
    .B(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__and2_1 _2264_ (.A(_0955_),
    .B(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__xor2_2 _2265_ (.A(_0955_),
    .B(_0957_),
    .X(_0959_));
 sky130_fd_sc_hd__a21oi_1 _2266_ (.A1(_0610_),
    .A2(_0780_),
    .B1(_0810_),
    .Y(_0960_));
 sky130_fd_sc_hd__and3_1 _2267_ (.A(_0913_),
    .B(_0916_),
    .C(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__a21oi_1 _2268_ (.A1(_0913_),
    .A2(_0916_),
    .B1(_0809_),
    .Y(_0962_));
 sky130_fd_sc_hd__a21oi_1 _2269_ (.A1(_0573_),
    .A2(_0610_),
    .B1(_0613_),
    .Y(_0963_));
 sky130_fd_sc_hd__a21o_1 _2270_ (.A1(_0573_),
    .A2(_0610_),
    .B1(_0613_),
    .X(_0964_));
 sky130_fd_sc_hd__o211a_1 _2271_ (.A1(_0717_),
    .A2(_0719_),
    .B1(_0963_),
    .C1(_0690_),
    .X(_0965_));
 sky130_fd_sc_hd__o211ai_1 _2272_ (.A1(_0717_),
    .A2(_0719_),
    .B1(_0964_),
    .C1(_0690_),
    .Y(_0966_));
 sky130_fd_sc_hd__o221a_1 _2273_ (.A1(_0612_),
    .A2(_0720_),
    .B1(_0961_),
    .B2(_0962_),
    .C1(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__a2111o_1 _2274_ (.A1(_0612_),
    .A2(_0721_),
    .B1(_0961_),
    .C1(_0962_),
    .D1(_0965_),
    .X(_0968_));
 sky130_fd_sc_hd__and2b_1 _2275_ (.A_N(_0967_),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__a21o_1 _2276_ (.A1(_0610_),
    .A2(_0968_),
    .B1(_0967_),
    .X(_0970_));
 sky130_fd_sc_hd__a21oi_1 _2277_ (.A1(_0959_),
    .A2(_0970_),
    .B1(_0958_),
    .Y(_0971_));
 sky130_fd_sc_hd__a211o_1 _2278_ (.A1(_0959_),
    .A2(_0970_),
    .B1(_0953_),
    .C1(_0958_),
    .X(_0972_));
 sky130_fd_sc_hd__nor2_1 _2279_ (.A(_0951_),
    .B(_0953_),
    .Y(_0973_));
 sky130_fd_sc_hd__nand2_1 _2280_ (.A(_0952_),
    .B(_0972_),
    .Y(_0974_));
 sky130_fd_sc_hd__a31o_1 _2281_ (.A1(_0945_),
    .A2(_0952_),
    .A3(_0972_),
    .B1(_0944_),
    .X(_0975_));
 sky130_fd_sc_hd__nand2_1 _2282_ (.A(_0936_),
    .B(_0938_),
    .Y(_0976_));
 sky130_fd_sc_hd__nand2b_1 _2283_ (.A_N(_0939_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__a21o_1 _2284_ (.A1(_0975_),
    .A2(_0976_),
    .B1(_0939_),
    .X(_0978_));
 sky130_fd_sc_hd__or2_1 _2285_ (.A(_0643_),
    .B(_0721_),
    .X(_0979_));
 sky130_fd_sc_hd__xnor2_1 _2286_ (.A(_0666_),
    .B(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__nor2_1 _2287_ (.A(_0839_),
    .B(_0917_),
    .Y(_0981_));
 sky130_fd_sc_hd__xnor2_1 _2288_ (.A(_0863_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__and2b_1 _2289_ (.A_N(_0980_),
    .B(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__xnor2_1 _2290_ (.A(_0980_),
    .B(_0982_),
    .Y(_0984_));
 sky130_fd_sc_hd__nor2_1 _2291_ (.A(_0724_),
    .B(_0921_),
    .Y(_0985_));
 sky130_fd_sc_hd__or2_1 _2292_ (.A(_0724_),
    .B(_0921_),
    .X(_0986_));
 sky130_fd_sc_hd__a211o_1 _2293_ (.A1(_0978_),
    .A2(_0984_),
    .B1(_0985_),
    .C1(_0983_),
    .X(_0987_));
 sky130_fd_sc_hd__a211oi_1 _2294_ (.A1(_0922_),
    .A2(_0987_),
    .B1(_0934_),
    .C1(_1166_),
    .Y(_0988_));
 sky130_fd_sc_hd__a211o_1 _2295_ (.A1(_0922_),
    .A2(_0987_),
    .B1(_0934_),
    .C1(_1166_),
    .X(_0989_));
 sky130_fd_sc_hd__o21a_1 _2296_ (.A1(net284),
    .A2(\gray_sobel0.sobel0.px_ready ),
    .B1(_0989_),
    .X(_0206_));
 sky130_fd_sc_hd__xor2_2 _2297_ (.A(_0610_),
    .B(_0969_),
    .X(_0990_));
 sky130_fd_sc_hd__o22a_1 _2298_ (.A1(net315),
    .A2(\gray_sobel0.sobel0.px_ready ),
    .B1(_0989_),
    .B2(_0990_),
    .X(_0207_));
 sky130_fd_sc_hd__xnor2_1 _2299_ (.A(_0959_),
    .B(_0970_),
    .Y(_0991_));
 sky130_fd_sc_hd__o2bb2a_1 _2300_ (.A1_N(_0988_),
    .A2_N(_0991_),
    .B1(net366),
    .B2(\gray_sobel0.sobel0.px_ready ),
    .X(_0208_));
 sky130_fd_sc_hd__xnor2_2 _2301_ (.A(_0971_),
    .B(_0973_),
    .Y(_0992_));
 sky130_fd_sc_hd__o22a_1 _2302_ (.A1(net292),
    .A2(\gray_sobel0.sobel0.px_ready ),
    .B1(_0989_),
    .B2(_0992_),
    .X(_0209_));
 sky130_fd_sc_hd__xnor2_1 _2303_ (.A(_0946_),
    .B(_0974_),
    .Y(_0993_));
 sky130_fd_sc_hd__o2bb2a_1 _2304_ (.A1_N(_0988_),
    .A2_N(_0993_),
    .B1(net319),
    .B2(\gray_sobel0.sobel0.px_ready ),
    .X(_0210_));
 sky130_fd_sc_hd__xnor2_1 _2305_ (.A(_0975_),
    .B(_0977_),
    .Y(_0994_));
 sky130_fd_sc_hd__o22a_1 _2306_ (.A1(net326),
    .A2(\gray_sobel0.sobel0.px_ready ),
    .B1(_0989_),
    .B2(_0994_),
    .X(_0211_));
 sky130_fd_sc_hd__xnor2_1 _2307_ (.A(_0978_),
    .B(_0984_),
    .Y(_0995_));
 sky130_fd_sc_hd__o2bb2a_1 _2308_ (.A1_N(_0988_),
    .A2_N(_0995_),
    .B1(net338),
    .B2(\gray_sobel0.sobel0.px_ready ),
    .X(_0212_));
 sky130_fd_sc_hd__a21o_1 _2309_ (.A1(_0922_),
    .A2(_0986_),
    .B1(_1166_),
    .X(_0996_));
 sky130_fd_sc_hd__o32a_1 _2310_ (.A1(_0934_),
    .A2(_0987_),
    .A3(_0996_),
    .B1(\gray_sobel0.sobel0.px_ready ),
    .B2(net277),
    .X(_0213_));
 sky130_fd_sc_hd__or4b_4 _2311_ (.A(\gray_sobel0.sobel0.counter_sobel[1] ),
    .B(\gray_sobel0.sobel0.counter_sobel[2] ),
    .C(\gray_sobel0.sobel0.counter_sobel[3] ),
    .D_N(\gray_sobel0.sobel0.counter_sobel[0] ),
    .X(_0997_));
 sky130_fd_sc_hd__nand2b_1 _2312_ (.A_N(\gray_sobel0.sobel0.counter_sobel[3] ),
    .B(\gray_sobel0.sobel0.counter_sobel[2] ),
    .Y(_0998_));
 sky130_fd_sc_hd__o21a_1 _2313_ (.A1(_0500_),
    .A2(_0998_),
    .B1(net33),
    .X(_0999_));
 sky130_fd_sc_hd__a211oi_4 _2314_ (.A1(net47),
    .A2(_0997_),
    .B1(_0999_),
    .C1(_1222_),
    .Y(_1000_));
 sky130_fd_sc_hd__mux2_1 _2315_ (.A0(net419),
    .A1(_0390_),
    .S(_1000_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2316_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[1] ),
    .A1(_0396_),
    .S(_1000_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2317_ (.A0(net393),
    .A1(_0402_),
    .S(_1000_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2318_ (.A0(net391),
    .A1(_0408_),
    .S(_1000_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2319_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[4] ),
    .A1(_0413_),
    .S(_1000_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[5] ),
    .A1(_0418_),
    .S(_1000_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2321_ (.A0(net358),
    .A1(_0423_),
    .S(_1000_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(net364),
    .A1(_0428_),
    .S(_1000_),
    .X(_0221_));
 sky130_fd_sc_hd__nor2_1 _2323_ (.A(_1219_),
    .B(_1221_),
    .Y(_1001_));
 sky130_fd_sc_hd__or2_1 _2324_ (.A(_1226_),
    .B(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__xnor2_1 _2325_ (.A(\gray_sobel0.sobel0.counter_sobel[0] ),
    .B(_1001_),
    .Y(_1003_));
 sky130_fd_sc_hd__and2_1 _2326_ (.A(net25),
    .B(_1003_),
    .X(_0222_));
 sky130_fd_sc_hd__a21o_1 _2327_ (.A1(net47),
    .A2(_1223_),
    .B1(\gray_sobel0.sobel0.next[0] ),
    .X(_1004_));
 sky130_fd_sc_hd__and3_1 _2328_ (.A(_1224_),
    .B(_0500_),
    .C(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _2329_ (.A0(_1005_),
    .A1(\gray_sobel0.sobel0.counter_sobel[1] ),
    .S(_1001_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _2330_ (.A(\gray_sobel0.sobel0.counter_sobel[1] ),
    .B(\gray_sobel0.sobel0.counter_sobel[0] ),
    .C(_1221_),
    .X(_1006_));
 sky130_fd_sc_hd__xnor2_1 _2331_ (.A(\gray_sobel0.sobel0.counter_sobel[2] ),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__nor2_1 _2332_ (.A(_1219_),
    .B(_1007_),
    .Y(_0224_));
 sky130_fd_sc_hd__or3b_1 _2333_ (.A(_1001_),
    .B(_0500_),
    .C_N(\gray_sobel0.sobel0.counter_sobel[2] ),
    .X(_1008_));
 sky130_fd_sc_hd__a211o_1 _2334_ (.A1(net33),
    .A2(_1225_),
    .B1(_1001_),
    .C1(net47),
    .X(_1009_));
 sky130_fd_sc_hd__xnor2_1 _2335_ (.A(\gray_sobel0.sobel0.counter_sobel[3] ),
    .B(_1008_),
    .Y(_1010_));
 sky130_fd_sc_hd__and2_1 _2336_ (.A(_1009_),
    .B(_1010_),
    .X(_0225_));
 sky130_fd_sc_hd__or3b_1 _2337_ (.A(\gray_sobel0.sobel0.counter_sobel[0] ),
    .B(_0998_),
    .C_N(\gray_sobel0.sobel0.counter_sobel[1] ),
    .X(_1011_));
 sky130_fd_sc_hd__a21oi_4 _2338_ (.A1(net33),
    .A2(_1011_),
    .B1(_0503_),
    .Y(_1012_));
 sky130_fd_sc_hd__mux2_1 _2339_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ),
    .A1(_0390_),
    .S(_1012_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2340_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ),
    .A1(_0396_),
    .S(_1012_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2341_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[2] ),
    .A1(_0402_),
    .S(_1012_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ),
    .A1(_0408_),
    .S(_1012_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ),
    .A1(_0413_),
    .S(_1012_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2344_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ),
    .A1(_0418_),
    .S(_1012_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2345_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[6] ),
    .A1(_0423_),
    .S(_1012_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ),
    .A1(_0428_),
    .S(_1012_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(net28),
    .A1(net25),
    .S(\gray_sobel0.sobel0.counter_pixels[0] ),
    .X(_0234_));
 sky130_fd_sc_hd__nand2_1 _2348_ (.A(\gray_sobel0.sobel0.counter_pixels[0] ),
    .B(\gray_sobel0.sobel0.counter_pixels[1] ),
    .Y(_1013_));
 sky130_fd_sc_hd__or2_1 _2349_ (.A(\gray_sobel0.sobel0.counter_pixels[0] ),
    .B(\gray_sobel0.sobel0.counter_pixels[1] ),
    .X(_1014_));
 sky130_fd_sc_hd__a32o_1 _2350_ (.A1(net28),
    .A2(_1013_),
    .A3(_1014_),
    .B1(net25),
    .B2(\gray_sobel0.sobel0.counter_pixels[1] ),
    .X(_0235_));
 sky130_fd_sc_hd__a21o_1 _2351_ (.A1(\gray_sobel0.sobel0.counter_pixels[0] ),
    .A2(\gray_sobel0.sobel0.counter_pixels[1] ),
    .B1(\gray_sobel0.sobel0.counter_pixels[2] ),
    .X(_1015_));
 sky130_fd_sc_hd__nand3_1 _2352_ (.A(\gray_sobel0.sobel0.counter_pixels[0] ),
    .B(\gray_sobel0.sobel0.counter_pixels[1] ),
    .C(\gray_sobel0.sobel0.counter_pixels[2] ),
    .Y(_1016_));
 sky130_fd_sc_hd__a32o_1 _2353_ (.A1(net28),
    .A2(_1015_),
    .A3(_1016_),
    .B1(net25),
    .B2(\gray_sobel0.sobel0.counter_pixels[2] ),
    .X(_0236_));
 sky130_fd_sc_hd__a31o_1 _2354_ (.A1(\gray_sobel0.sobel0.counter_pixels[0] ),
    .A2(\gray_sobel0.sobel0.counter_pixels[1] ),
    .A3(\gray_sobel0.sobel0.counter_pixels[2] ),
    .B1(\gray_sobel0.sobel0.counter_pixels[3] ),
    .X(_1017_));
 sky130_fd_sc_hd__and4_1 _2355_ (.A(\gray_sobel0.sobel0.counter_pixels[0] ),
    .B(\gray_sobel0.sobel0.counter_pixels[1] ),
    .C(\gray_sobel0.sobel0.counter_pixels[3] ),
    .D(\gray_sobel0.sobel0.counter_pixels[2] ),
    .X(_1018_));
 sky130_fd_sc_hd__inv_2 _2356_ (.A(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__a32o_1 _2357_ (.A1(net28),
    .A2(_1017_),
    .A3(_1019_),
    .B1(net25),
    .B2(net390),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _2358_ (.A(\gray_sobel0.sobel0.counter_pixels[4] ),
    .B(_1018_),
    .X(_1020_));
 sky130_fd_sc_hd__nand2_1 _2359_ (.A(\gray_sobel0.sobel0.counter_pixels[4] ),
    .B(_1018_),
    .Y(_1021_));
 sky130_fd_sc_hd__a32o_1 _2360_ (.A1(net26),
    .A2(_1020_),
    .A3(_1021_),
    .B1(net25),
    .B2(\gray_sobel0.sobel0.counter_pixels[4] ),
    .X(_0238_));
 sky130_fd_sc_hd__a21o_1 _2361_ (.A1(\gray_sobel0.sobel0.counter_pixels[4] ),
    .A2(_1018_),
    .B1(\gray_sobel0.sobel0.counter_pixels[5] ),
    .X(_1022_));
 sky130_fd_sc_hd__and3_1 _2362_ (.A(\gray_sobel0.sobel0.counter_pixels[5] ),
    .B(\gray_sobel0.sobel0.counter_pixels[4] ),
    .C(_1018_),
    .X(_1023_));
 sky130_fd_sc_hd__inv_2 _2363_ (.A(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__a32o_1 _2364_ (.A1(net26),
    .A2(_1022_),
    .A3(_1024_),
    .B1(net25),
    .B2(net374),
    .X(_0239_));
 sky130_fd_sc_hd__or2_1 _2365_ (.A(\gray_sobel0.sobel0.counter_pixels[6] ),
    .B(_1023_),
    .X(_1025_));
 sky130_fd_sc_hd__and2_1 _2366_ (.A(\gray_sobel0.sobel0.counter_pixels[6] ),
    .B(_1023_),
    .X(_1026_));
 sky130_fd_sc_hd__inv_2 _2367_ (.A(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__a32o_1 _2368_ (.A1(net26),
    .A2(_1025_),
    .A3(_1027_),
    .B1(net25),
    .B2(net408),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _2369_ (.A(\gray_sobel0.sobel0.counter_pixels[7] ),
    .B(_1026_),
    .X(_1028_));
 sky130_fd_sc_hd__nand2_1 _2370_ (.A(\gray_sobel0.sobel0.counter_pixels[7] ),
    .B(_1026_),
    .Y(_1029_));
 sky130_fd_sc_hd__a32o_1 _2371_ (.A1(net26),
    .A2(_1028_),
    .A3(_1029_),
    .B1(net25),
    .B2(\gray_sobel0.sobel0.counter_pixels[7] ),
    .X(_0241_));
 sky130_fd_sc_hd__a31o_1 _2372_ (.A1(\gray_sobel0.sobel0.counter_pixels[7] ),
    .A2(\gray_sobel0.sobel0.counter_pixels[6] ),
    .A3(_1023_),
    .B1(\gray_sobel0.sobel0.counter_pixels[8] ),
    .X(_1030_));
 sky130_fd_sc_hd__and3_1 _2373_ (.A(\gray_sobel0.sobel0.counter_pixels[7] ),
    .B(\gray_sobel0.sobel0.counter_pixels[8] ),
    .C(_1026_),
    .X(_1031_));
 sky130_fd_sc_hd__inv_2 _2374_ (.A(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__a32o_1 _2375_ (.A1(net26),
    .A2(_1030_),
    .A3(_1032_),
    .B1(net24),
    .B2(net399),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _2376_ (.A(\gray_sobel0.sobel0.counter_pixels[9] ),
    .B(_1031_),
    .X(_1033_));
 sky130_fd_sc_hd__nand2_1 _2377_ (.A(\gray_sobel0.sobel0.counter_pixels[9] ),
    .B(_1031_),
    .Y(_1034_));
 sky130_fd_sc_hd__a32o_1 _2378_ (.A1(net26),
    .A2(_1033_),
    .A3(_1034_),
    .B1(net24),
    .B2(net459),
    .X(_0243_));
 sky130_fd_sc_hd__and3_1 _2379_ (.A(\gray_sobel0.sobel0.counter_pixels[9] ),
    .B(\gray_sobel0.sobel0.counter_pixels[10] ),
    .C(_1031_),
    .X(_1035_));
 sky130_fd_sc_hd__a21oi_1 _2380_ (.A1(\gray_sobel0.sobel0.counter_pixels[9] ),
    .A2(_1031_),
    .B1(\gray_sobel0.sobel0.counter_pixels[10] ),
    .Y(_1036_));
 sky130_fd_sc_hd__nor2_1 _2381_ (.A(_1035_),
    .B(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__a22o_1 _2382_ (.A1(net446),
    .A2(net24),
    .B1(_1037_),
    .B2(net28),
    .X(_0244_));
 sky130_fd_sc_hd__and2_1 _2383_ (.A(\gray_sobel0.sobel0.counter_pixels[11] ),
    .B(_1035_),
    .X(_1038_));
 sky130_fd_sc_hd__o21ai_1 _2384_ (.A1(\gray_sobel0.sobel0.counter_pixels[11] ),
    .A2(_1035_),
    .B1(net28),
    .Y(_1039_));
 sky130_fd_sc_hd__a2bb2o_1 _2385_ (.A1_N(_1038_),
    .A2_N(_1039_),
    .B1(\gray_sobel0.sobel0.counter_pixels[11] ),
    .B2(net24),
    .X(_0245_));
 sky130_fd_sc_hd__and3_1 _2386_ (.A(\gray_sobel0.sobel0.counter_pixels[11] ),
    .B(\gray_sobel0.sobel0.counter_pixels[12] ),
    .C(_1035_),
    .X(_1040_));
 sky130_fd_sc_hd__o21ai_1 _2387_ (.A1(\gray_sobel0.sobel0.counter_pixels[12] ),
    .A2(_1038_),
    .B1(net27),
    .Y(_1041_));
 sky130_fd_sc_hd__a2bb2o_1 _2388_ (.A1_N(_1040_),
    .A2_N(_1041_),
    .B1(net435),
    .B2(net24),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_1 _2389_ (.A(\gray_sobel0.sobel0.counter_pixels[13] ),
    .B(_1040_),
    .Y(_1042_));
 sky130_fd_sc_hd__or2_1 _2390_ (.A(\gray_sobel0.sobel0.counter_pixels[13] ),
    .B(_1040_),
    .X(_1043_));
 sky130_fd_sc_hd__a32o_1 _2391_ (.A1(net27),
    .A2(_1042_),
    .A3(_1043_),
    .B1(net23),
    .B2(\gray_sobel0.sobel0.counter_pixels[13] ),
    .X(_0247_));
 sky130_fd_sc_hd__and3_1 _2392_ (.A(\gray_sobel0.sobel0.counter_pixels[13] ),
    .B(\gray_sobel0.sobel0.counter_pixels[14] ),
    .C(_1040_),
    .X(_1044_));
 sky130_fd_sc_hd__inv_2 _2393_ (.A(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a21o_1 _2394_ (.A1(\gray_sobel0.sobel0.counter_pixels[13] ),
    .A2(_1040_),
    .B1(\gray_sobel0.sobel0.counter_pixels[14] ),
    .X(_1046_));
 sky130_fd_sc_hd__a32o_1 _2395_ (.A1(net26),
    .A2(_1045_),
    .A3(_1046_),
    .B1(net23),
    .B2(net379),
    .X(_0248_));
 sky130_fd_sc_hd__and2_1 _2396_ (.A(\gray_sobel0.sobel0.counter_pixels[15] ),
    .B(_1044_),
    .X(_1047_));
 sky130_fd_sc_hd__o21ai_1 _2397_ (.A1(\gray_sobel0.sobel0.counter_pixels[15] ),
    .A2(_1044_),
    .B1(net26),
    .Y(_1048_));
 sky130_fd_sc_hd__a2bb2o_1 _2398_ (.A1_N(_1047_),
    .A2_N(_1048_),
    .B1(\gray_sobel0.sobel0.counter_pixels[15] ),
    .B2(net23),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _2399_ (.A(\gray_sobel0.sobel0.counter_pixels[16] ),
    .B(_1047_),
    .Y(_1049_));
 sky130_fd_sc_hd__or2_1 _2400_ (.A(\gray_sobel0.sobel0.counter_pixels[16] ),
    .B(_1047_),
    .X(_1050_));
 sky130_fd_sc_hd__a32o_1 _2401_ (.A1(net26),
    .A2(_1049_),
    .A3(_1050_),
    .B1(net23),
    .B2(\gray_sobel0.sobel0.counter_pixels[16] ),
    .X(_0250_));
 sky130_fd_sc_hd__and3_1 _2402_ (.A(\gray_sobel0.sobel0.counter_pixels[17] ),
    .B(\gray_sobel0.sobel0.counter_pixels[16] ),
    .C(_1047_),
    .X(_1051_));
 sky130_fd_sc_hd__inv_2 _2403_ (.A(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__a31o_1 _2404_ (.A1(\gray_sobel0.sobel0.counter_pixels[15] ),
    .A2(\gray_sobel0.sobel0.counter_pixels[16] ),
    .A3(_1044_),
    .B1(\gray_sobel0.sobel0.counter_pixels[17] ),
    .X(_1053_));
 sky130_fd_sc_hd__a32o_1 _2405_ (.A1(net26),
    .A2(_1052_),
    .A3(_1053_),
    .B1(net23),
    .B2(net372),
    .X(_0251_));
 sky130_fd_sc_hd__and2_1 _2406_ (.A(\gray_sobel0.sobel0.counter_pixels[18] ),
    .B(_1051_),
    .X(_1054_));
 sky130_fd_sc_hd__o21ai_1 _2407_ (.A1(\gray_sobel0.sobel0.counter_pixels[18] ),
    .A2(_1051_),
    .B1(net27),
    .Y(_1055_));
 sky130_fd_sc_hd__a2bb2o_1 _2408_ (.A1_N(_1054_),
    .A2_N(_1055_),
    .B1(\gray_sobel0.sobel0.counter_pixels[18] ),
    .B2(net23),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _2409_ (.A(\gray_sobel0.sobel0.counter_pixels[19] ),
    .B(_1054_),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_1 _2410_ (.A(\gray_sobel0.sobel0.counter_pixels[19] ),
    .B(_1054_),
    .Y(_1057_));
 sky130_fd_sc_hd__a32o_1 _2411_ (.A1(net27),
    .A2(_1056_),
    .A3(_1057_),
    .B1(net23),
    .B2(\gray_sobel0.sobel0.counter_pixels[19] ),
    .X(_0253_));
 sky130_fd_sc_hd__a31o_1 _2412_ (.A1(\gray_sobel0.sobel0.counter_pixels[19] ),
    .A2(\gray_sobel0.sobel0.counter_pixels[18] ),
    .A3(_1051_),
    .B1(\gray_sobel0.sobel0.counter_pixels[20] ),
    .X(_1058_));
 sky130_fd_sc_hd__and3_1 _2413_ (.A(\gray_sobel0.sobel0.counter_pixels[19] ),
    .B(\gray_sobel0.sobel0.counter_pixels[20] ),
    .C(_1054_),
    .X(_1059_));
 sky130_fd_sc_hd__inv_2 _2414_ (.A(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__a32o_1 _2415_ (.A1(net27),
    .A2(_1058_),
    .A3(_1060_),
    .B1(net23),
    .B2(net402),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _2416_ (.A(\gray_sobel0.sobel0.counter_pixels[21] ),
    .B(_1059_),
    .Y(_1061_));
 sky130_fd_sc_hd__or2_1 _2417_ (.A(\gray_sobel0.sobel0.counter_pixels[21] ),
    .B(_1059_),
    .X(_1062_));
 sky130_fd_sc_hd__a32o_1 _2418_ (.A1(net27),
    .A2(_1061_),
    .A3(_1062_),
    .B1(net23),
    .B2(\gray_sobel0.sobel0.counter_pixels[21] ),
    .X(_0255_));
 sky130_fd_sc_hd__nand3_1 _2419_ (.A(\gray_sobel0.sobel0.counter_pixels[21] ),
    .B(\gray_sobel0.sobel0.counter_pixels[22] ),
    .C(_1059_),
    .Y(_1063_));
 sky130_fd_sc_hd__a21o_1 _2420_ (.A1(net27),
    .A2(_1063_),
    .B1(net23),
    .X(_1064_));
 sky130_fd_sc_hd__a31o_1 _2421_ (.A1(\gray_sobel0.sobel0.counter_pixels[21] ),
    .A2(net27),
    .A3(_1059_),
    .B1(\gray_sobel0.sobel0.counter_pixels[22] ),
    .X(_1065_));
 sky130_fd_sc_hd__and2_1 _2422_ (.A(_1064_),
    .B(_1065_),
    .X(_0256_));
 sky130_fd_sc_hd__or3b_1 _2423_ (.A(_1063_),
    .B(\gray_sobel0.sobel0.counter_pixels[23] ),
    .C_N(net27),
    .X(_1066_));
 sky130_fd_sc_hd__a21bo_1 _2424_ (.A1(net297),
    .A2(_1064_),
    .B1_N(_1066_),
    .X(_0257_));
 sky130_fd_sc_hd__a21o_1 _2425_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[0] ),
    .A2(net43),
    .B1(_0505_),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(_1067_),
    .A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[0] ),
    .S(_0502_),
    .X(_0258_));
 sky130_fd_sc_hd__a21o_1 _2427_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[1] ),
    .A2(net43),
    .B1(_0507_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _2428_ (.A0(_1068_),
    .A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[1] ),
    .S(_0502_),
    .X(_0259_));
 sky130_fd_sc_hd__a21o_1 _2429_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[2] ),
    .A2(net45),
    .B1(_0509_),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _2430_ (.A0(_1069_),
    .A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[2] ),
    .S(_0502_),
    .X(_0260_));
 sky130_fd_sc_hd__a21o_1 _2431_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[3] ),
    .A2(net44),
    .B1(_0511_),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _2432_ (.A0(_1070_),
    .A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[3] ),
    .S(_0502_),
    .X(_0261_));
 sky130_fd_sc_hd__a21o_1 _2433_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[4] ),
    .A2(net45),
    .B1(_0513_),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(_1071_),
    .A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[4] ),
    .S(_0502_),
    .X(_0262_));
 sky130_fd_sc_hd__a21o_1 _2435_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[5] ),
    .A2(net46),
    .B1(_0515_),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(_1072_),
    .A1(net453),
    .S(_0502_),
    .X(_0263_));
 sky130_fd_sc_hd__a21o_1 _2437_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[6] ),
    .A2(net48),
    .B1(_0517_),
    .X(_1073_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(_1073_),
    .A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[6] ),
    .S(_0502_),
    .X(_0264_));
 sky130_fd_sc_hd__a21o_1 _2439_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[7] ),
    .A2(net47),
    .B1(_0519_),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(_1074_),
    .A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[7] ),
    .S(_0502_),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_4 _2441_ (.A1(net33),
    .A2(_0997_),
    .B1(_0503_),
    .Y(_1075_));
 sky130_fd_sc_hd__a21o_1 _2442_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[0] ),
    .A2(net42),
    .B1(_0505_),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_1 _2443_ (.A0(net245),
    .A1(_1076_),
    .S(_1075_),
    .X(_0266_));
 sky130_fd_sc_hd__a21o_1 _2444_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[1] ),
    .A2(net42),
    .B1(_0507_),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(net249),
    .A1(_1077_),
    .S(_1075_),
    .X(_0267_));
 sky130_fd_sc_hd__a21o_1 _2446_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[2] ),
    .A2(net43),
    .B1(_0509_),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(net248),
    .A1(_1078_),
    .S(_1075_),
    .X(_0268_));
 sky130_fd_sc_hd__a21o_1 _2448_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[3] ),
    .A2(net44),
    .B1(_0511_),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _2449_ (.A0(net241),
    .A1(_1079_),
    .S(_1075_),
    .X(_0269_));
 sky130_fd_sc_hd__a21o_1 _2450_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[4] ),
    .A2(net45),
    .B1(_0513_),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_1 _2451_ (.A0(net202),
    .A1(_1080_),
    .S(_1075_),
    .X(_0270_));
 sky130_fd_sc_hd__a21o_1 _2452_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[5] ),
    .A2(net46),
    .B1(_0515_),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[5] ),
    .A1(_1081_),
    .S(_1075_),
    .X(_0271_));
 sky130_fd_sc_hd__a21o_1 _2454_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[6] ),
    .A2(net46),
    .B1(_0517_),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(net240),
    .A1(_1082_),
    .S(_1075_),
    .X(_0272_));
 sky130_fd_sc_hd__a21o_1 _2456_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[7] ),
    .A2(net48),
    .B1(_0519_),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _2457_ (.A0(net234),
    .A1(_1083_),
    .S(_1075_),
    .X(_0273_));
 sky130_fd_sc_hd__or3b_1 _2458_ (.A(_0998_),
    .B(\gray_sobel0.sobel0.counter_sobel[1] ),
    .C_N(\gray_sobel0.sobel0.counter_sobel[0] ),
    .X(_1084_));
 sky130_fd_sc_hd__a21oi_4 _2459_ (.A1(net33),
    .A2(_1084_),
    .B1(_0503_),
    .Y(_1085_));
 sky130_fd_sc_hd__a21o_1 _2460_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ),
    .A2(net42),
    .B1(_0505_),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _2461_ (.A0(net247),
    .A1(_1086_),
    .S(_1085_),
    .X(_0274_));
 sky130_fd_sc_hd__a21o_1 _2462_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ),
    .A2(net42),
    .B1(_0507_),
    .X(_1087_));
 sky130_fd_sc_hd__mux2_1 _2463_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[1] ),
    .A1(_1087_),
    .S(_1085_),
    .X(_0275_));
 sky130_fd_sc_hd__a21o_1 _2464_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ),
    .A2(net43),
    .B1(_0509_),
    .X(_1088_));
 sky130_fd_sc_hd__mux2_1 _2465_ (.A0(net244),
    .A1(_1088_),
    .S(_1085_),
    .X(_0276_));
 sky130_fd_sc_hd__a21o_1 _2466_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ),
    .A2(net44),
    .B1(_0511_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(net243),
    .A1(_1089_),
    .S(_1085_),
    .X(_0277_));
 sky130_fd_sc_hd__a21o_1 _2468_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ),
    .A2(net44),
    .B1(_0513_),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[4] ),
    .A1(_1090_),
    .S(_1085_),
    .X(_0278_));
 sky130_fd_sc_hd__a21o_1 _2470_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[5] ),
    .A2(net46),
    .B1(_0515_),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_1 _2471_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[5] ),
    .A1(_1091_),
    .S(_1085_),
    .X(_0279_));
 sky130_fd_sc_hd__a21o_1 _2472_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ),
    .A2(net49),
    .B1(_0517_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_1 _2473_ (.A0(net203),
    .A1(_1092_),
    .S(_1085_),
    .X(_0280_));
 sky130_fd_sc_hd__a21o_1 _2474_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ),
    .A2(net48),
    .B1(_0519_),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _2475_ (.A0(net237),
    .A1(_1093_),
    .S(_1085_),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_4 _2476_ (.A1(\gray_sobel0.sobel0.next[0] ),
    .A2(_1223_),
    .B1(_0503_),
    .Y(_1094_));
 sky130_fd_sc_hd__a21o_1 _2477_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[0] ),
    .A2(net42),
    .B1(_0505_),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[0] ),
    .A1(_1095_),
    .S(_1094_),
    .X(_0282_));
 sky130_fd_sc_hd__a21o_1 _2479_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[1] ),
    .A2(net43),
    .B1(_0507_),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _2480_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[1] ),
    .A1(_1096_),
    .S(_1094_),
    .X(_0283_));
 sky130_fd_sc_hd__a21o_1 _2481_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[2] ),
    .A2(net43),
    .B1(_0509_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[2] ),
    .A1(_1097_),
    .S(_1094_),
    .X(_0284_));
 sky130_fd_sc_hd__a21o_1 _2483_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[3] ),
    .A2(net44),
    .B1(_0511_),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _2484_ (.A0(net199),
    .A1(_1098_),
    .S(_1094_),
    .X(_0285_));
 sky130_fd_sc_hd__a21o_1 _2485_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[4] ),
    .A2(net45),
    .B1(_0513_),
    .X(_1099_));
 sky130_fd_sc_hd__mux2_1 _2486_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[4] ),
    .A1(_1099_),
    .S(_1094_),
    .X(_0286_));
 sky130_fd_sc_hd__a21o_1 _2487_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[5] ),
    .A2(net46),
    .B1(_0515_),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _2488_ (.A0(net198),
    .A1(_1100_),
    .S(_1094_),
    .X(_0287_));
 sky130_fd_sc_hd__a21o_1 _2489_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[6] ),
    .A2(net46),
    .B1(_0517_),
    .X(_1101_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[6] ),
    .A1(_1101_),
    .S(_1094_),
    .X(_0288_));
 sky130_fd_sc_hd__a21o_1 _2491_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[7] ),
    .A2(net47),
    .B1(_0519_),
    .X(_1102_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[7] ),
    .A1(_1102_),
    .S(_1094_),
    .X(_0289_));
 sky130_fd_sc_hd__o21a_1 _2493_ (.A1(_1224_),
    .A2(_0998_),
    .B1(net33),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_4 _2494_ (.A(_0503_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__a21o_1 _2495_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[0] ),
    .A2(net42),
    .B1(_0505_),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(net291),
    .A1(_1105_),
    .S(_1104_),
    .X(_0290_));
 sky130_fd_sc_hd__a21o_1 _2497_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[1] ),
    .A2(net42),
    .B1(_0507_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(net281),
    .A1(_1106_),
    .S(_1104_),
    .X(_0291_));
 sky130_fd_sc_hd__a21o_1 _2499_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[2] ),
    .A2(net43),
    .B1(_0509_),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_1 _2500_ (.A0(net283),
    .A1(_1107_),
    .S(_1104_),
    .X(_0292_));
 sky130_fd_sc_hd__a21o_1 _2501_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[3] ),
    .A2(net44),
    .B1(_0511_),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(net288),
    .A1(_1108_),
    .S(_1104_),
    .X(_0293_));
 sky130_fd_sc_hd__a21o_1 _2503_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[4] ),
    .A2(net44),
    .B1(_0513_),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(net285),
    .A1(_1109_),
    .S(_1104_),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _2505_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[5] ),
    .A2(net46),
    .B1(_0515_),
    .X(_1110_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(net286),
    .A1(_1110_),
    .S(_1104_),
    .X(_0295_));
 sky130_fd_sc_hd__a21o_1 _2507_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[6] ),
    .A2(net46),
    .B1(_0517_),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(net314),
    .A1(_1111_),
    .S(_1104_),
    .X(_0296_));
 sky130_fd_sc_hd__a21o_1 _2509_ (.A1(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[7] ),
    .A2(net48),
    .B1(_0519_),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(net293),
    .A1(_1112_),
    .S(_1104_),
    .X(_0297_));
 sky130_fd_sc_hd__xnor2_1 _2511_ (.A(\lfsr0.lfsr_out[3] ),
    .B(\lfsr0.lfsr_out[12] ),
    .Y(_1113_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(\lfsr0.seed_reg[0] ),
    .A1(_1113_),
    .S(net66),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _2513_ (.A0(\lfsr0.lfsr_out[0] ),
    .A1(_1114_),
    .S(net30),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(\lfsr0.seed_reg[1] ),
    .A1(\lfsr0.lfsr_out[0] ),
    .S(net66),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _2515_ (.A0(\lfsr0.lfsr_out[1] ),
    .A1(_1115_),
    .S(net30),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(\lfsr0.seed_reg[2] ),
    .A1(\lfsr0.lfsr_out[1] ),
    .S(net66),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(\lfsr0.lfsr_out[2] ),
    .A1(_1116_),
    .S(net30),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(\lfsr0.seed_reg[3] ),
    .A1(\lfsr0.lfsr_out[2] ),
    .S(net66),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(\lfsr0.lfsr_out[3] ),
    .A1(_1117_),
    .S(net30),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(\lfsr0.seed_reg[4] ),
    .A1(\lfsr0.lfsr_out[3] ),
    .S(net67),
    .X(_1118_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(\lfsr0.lfsr_out[4] ),
    .A1(_1118_),
    .S(net31),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(\lfsr0.seed_reg[5] ),
    .A1(\lfsr0.lfsr_out[4] ),
    .S(net67),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(\lfsr0.lfsr_out[5] ),
    .A1(_1119_),
    .S(net31),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(\lfsr0.seed_reg[6] ),
    .A1(\lfsr0.lfsr_out[5] ),
    .S(net68),
    .X(_1120_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(\lfsr0.lfsr_out[6] ),
    .A1(_1120_),
    .S(net32),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\lfsr0.seed_reg[7] ),
    .A1(\lfsr0.lfsr_out[6] ),
    .S(net68),
    .X(_1121_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(\lfsr0.lfsr_out[7] ),
    .A1(_1121_),
    .S(net32),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(\lfsr0.seed_reg[8] ),
    .A1(\lfsr0.lfsr_out[7] ),
    .S(net68),
    .X(_1122_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(\lfsr0.lfsr_out[8] ),
    .A1(_1122_),
    .S(net32),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(\lfsr0.seed_reg[9] ),
    .A1(\lfsr0.lfsr_out[8] ),
    .S(net67),
    .X(_1123_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(\lfsr0.lfsr_out[9] ),
    .A1(_1123_),
    .S(net31),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(\lfsr0.seed_reg[10] ),
    .A1(\lfsr0.lfsr_out[9] ),
    .S(net66),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(\lfsr0.lfsr_out[10] ),
    .A1(_1124_),
    .S(net30),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(\lfsr0.seed_reg[11] ),
    .A1(\lfsr0.lfsr_out[10] ),
    .S(net66),
    .X(_1125_));
 sky130_fd_sc_hd__mux2_1 _2535_ (.A0(\lfsr0.lfsr_out[11] ),
    .A1(_1125_),
    .S(net30),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(\lfsr0.seed_reg[12] ),
    .A1(\lfsr0.lfsr_out[11] ),
    .S(net66),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(\lfsr0.lfsr_out[12] ),
    .A1(_1126_),
    .S(net30),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(\lfsr0.seed_reg[13] ),
    .A1(\lfsr0.lfsr_out[12] ),
    .S(net66),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(\lfsr0.lfsr_out[13] ),
    .A1(_1127_),
    .S(net30),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(\lfsr0.seed_reg[14] ),
    .A1(\lfsr0.lfsr_out[13] ),
    .S(net66),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(\lfsr0.lfsr_out[14] ),
    .A1(_1128_),
    .S(net30),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(\lfsr0.seed_reg[15] ),
    .A1(\lfsr0.lfsr_out[14] ),
    .S(net67),
    .X(_1129_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(\lfsr0.lfsr_out[15] ),
    .A1(_1129_),
    .S(net31),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(\lfsr0.seed_reg[16] ),
    .A1(\lfsr0.lfsr_out[15] ),
    .S(net68),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(\lfsr0.lfsr_out[16] ),
    .A1(_1130_),
    .S(net32),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(\lfsr0.seed_reg[17] ),
    .A1(\lfsr0.lfsr_out[16] ),
    .S(net68),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_1 _2547_ (.A0(\lfsr0.lfsr_out[17] ),
    .A1(_1131_),
    .S(net32),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(\lfsr0.seed_reg[18] ),
    .A1(\lfsr0.lfsr_out[17] ),
    .S(net68),
    .X(_1132_));
 sky130_fd_sc_hd__mux2_1 _2549_ (.A0(\lfsr0.lfsr_out[18] ),
    .A1(_1132_),
    .S(net32),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(\lfsr0.seed_reg[19] ),
    .A1(\lfsr0.lfsr_out[18] ),
    .S(net68),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(\lfsr0.lfsr_out[19] ),
    .A1(_1133_),
    .S(net32),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(\lfsr0.seed_reg[20] ),
    .A1(\lfsr0.lfsr_out[19] ),
    .S(net67),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(\lfsr0.lfsr_out[20] ),
    .A1(_1134_),
    .S(net31),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(\lfsr0.seed_reg[21] ),
    .A1(\lfsr0.lfsr_out[20] ),
    .S(net67),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(\lfsr0.lfsr_out[21] ),
    .A1(_1135_),
    .S(net31),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2556_ (.A0(\lfsr0.seed_reg[22] ),
    .A1(\lfsr0.lfsr_out[21] ),
    .S(net66),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(\lfsr0.lfsr_out[22] ),
    .A1(_1136_),
    .S(net30),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(\lfsr0.seed_reg[23] ),
    .A1(\lfsr0.lfsr_out[22] ),
    .S(net67),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(\lfsr0.lfsr_out[23] ),
    .A1(_1137_),
    .S(net31),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ),
    .A1(_0390_),
    .S(net29),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ),
    .A1(_0396_),
    .S(net29),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ),
    .A1(_0402_),
    .S(net29),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ),
    .A1(_0408_),
    .S(net29),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _2564_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ),
    .A1(_0413_),
    .S(net29),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(net438),
    .A1(_0418_),
    .S(net29),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ),
    .A1(_0423_),
    .S(net29),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ),
    .A1(_0428_),
    .S(net29),
    .X(_0329_));
 sky130_fd_sc_hd__and2b_1 _2568_ (.A_N(net71),
    .B(in_lfsr_rdy),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(net327),
    .A1(\input_data[0] ),
    .S(net55),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(net324),
    .A1(\input_data[1] ),
    .S(net54),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(net350),
    .A1(\input_data[2] ),
    .S(net55),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(net375),
    .A1(\input_data[3] ),
    .S(net54),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(net352),
    .A1(\input_data[4] ),
    .S(net55),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(net332),
    .A1(\input_data[5] ),
    .S(net55),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(net328),
    .A1(\input_data[6] ),
    .S(net55),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(net367),
    .A1(\input_data[7] ),
    .S(net55),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _2577_ (.A0(net348),
    .A1(\input_data[8] ),
    .S(net56),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(net343),
    .A1(\input_data[9] ),
    .S(net56),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(net321),
    .A1(\input_data[10] ),
    .S(net54),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(net349),
    .A1(\input_data[11] ),
    .S(net55),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _2581_ (.A0(net331),
    .A1(\input_data[12] ),
    .S(net54),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(net336),
    .A1(\input_data[13] ),
    .S(net54),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(net354),
    .A1(\input_data[14] ),
    .S(net54),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(net320),
    .A1(\input_data[15] ),
    .S(net54),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(net368),
    .A1(\input_data[16] ),
    .S(net55),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(net341),
    .A1(\input_data[17] ),
    .S(net55),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(net339),
    .A1(\input_data[18] ),
    .S(net56),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(net356),
    .A1(\input_data[19] ),
    .S(net56),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(net322),
    .A1(\input_data[20] ),
    .S(net56),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(net362),
    .A1(\input_data[21] ),
    .S(net54),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(net344),
    .A1(\input_data[22] ),
    .S(net54),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(net346),
    .A1(\input_data[23] ),
    .S(net54),
    .X(_0353_));
 sky130_fd_sc_hd__and3_1 _2593_ (.A(in_data_rdy),
    .B(net74),
    .C(\lfsr0.config_i ),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _2594_ (.A0(\lfsr0.stop_reg[0] ),
    .A1(\input_data[0] ),
    .S(net57),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(net397),
    .A1(\input_data[1] ),
    .S(net57),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(net417),
    .A1(\input_data[2] ),
    .S(net59),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(\lfsr0.stop_reg[3] ),
    .A1(net411),
    .S(net57),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(\lfsr0.stop_reg[4] ),
    .A1(net394),
    .S(net58),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(net448),
    .A1(\input_data[5] ),
    .S(net58),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(net450),
    .A1(\input_data[6] ),
    .S(net58),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(net431),
    .A1(\input_data[7] ),
    .S(net58),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(net436),
    .A1(\input_data[8] ),
    .S(net58),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(net447),
    .A1(\input_data[9] ),
    .S(net59),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(net454),
    .A1(\input_data[10] ),
    .S(net57),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _2605_ (.A0(net455),
    .A1(\input_data[11] ),
    .S(net59),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _2606_ (.A0(net422),
    .A1(\input_data[12] ),
    .S(net57),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(net420),
    .A1(\input_data[13] ),
    .S(net57),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _2608_ (.A0(\lfsr0.stop_reg[14] ),
    .A1(net433),
    .S(net57),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(net457),
    .A1(\input_data[15] ),
    .S(net57),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(\lfsr0.stop_reg[16] ),
    .A1(net412),
    .S(net59),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(net443),
    .A1(net442),
    .S(net58),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(net439),
    .A1(net437),
    .S(net58),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(net445),
    .A1(net432),
    .S(net58),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _2614_ (.A0(net424),
    .A1(\input_data[20] ),
    .S(net58),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(\lfsr0.stop_reg[21] ),
    .A1(net444),
    .S(net57),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _2616_ (.A0(net414),
    .A1(\input_data[22] ),
    .S(net57),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(net426),
    .A1(\input_data[23] ),
    .S(net58),
    .X(_0377_));
 sky130_fd_sc_hd__inv_2 _2618_ (.A(net120),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _2619_ (.A(net120),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _2620_ (.A(net120),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _2621_ (.A(net123),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _2622_ (.A(net123),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _2623_ (.A(net120),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _2624_ (.A(net120),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _2625_ (.A(net120),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _2626_ (.A(net120),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _2627_ (.A(net120),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _2628_ (.A(net120),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _2629_ (.A(net120),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _2630_ (.A(net121),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _2631_ (.A(net121),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _2632_ (.A(net121),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _2633_ (.A(net118),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _2634_ (.A(net118),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _2635_ (.A(net118),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _2636_ (.A(net118),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _2637_ (.A(net118),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _2638_ (.A(net118),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _2639_ (.A(net118),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _2640_ (.A(net118),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _2641_ (.A(net119),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _2642_ (.A(net119),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _2643_ (.A(net119),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _2644_ (.A(net119),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _2645_ (.A(net118),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _2646_ (.A(net119),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _2648__3 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _2649__4 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _2650__5 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _2651__6 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _2653__7 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _2652_ (.A(net118),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _2654__8 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _2655__9 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _2656__10 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _2657__11 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _2658__12 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _2659__13 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _2660__14 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _2661__15 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _2662__16 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _2663__17 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _2664__18 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _2665__19 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _2666__20 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _2667__21 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _2668__22 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _2669__23 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _2670__24 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _2671__25 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _2672__26 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _2673__27 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _2674__28 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _2675__29 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _2676__30 (.A(clknet_2_3__leaf_ui_in[1]),
    .Y(net170));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__inv_2 _2677_ (.A(net123),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _2678_ (.A(net122),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _2679_ (.A(net122),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _2680_ (.A(net122),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _2681_ (.A(net122),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _2682_ (.A(net116),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _2683_ (.A(net115),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _2684_ (.A(net116),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _2685_ (.A(net116),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _2686_ (.A(net116),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _2687_ (.A(net115),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _2688_ (.A(net115),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _2689_ (.A(net115),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _2690_ (.A(net115),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _2691_ (.A(net115),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _2692_ (.A(net115),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _2693_ (.A(net115),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _2694_ (.A(net115),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _2695_ (.A(net115),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _2696_ (.A(net117),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _2697_ (.A(net117),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _2698_ (.A(net117),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _2699_ (.A(net116),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _2700_ (.A(net117),
    .Y(_0125_));
 sky130_fd_sc_hd__dfxtp_2 _2701_ (.CLK(clknet_leaf_11_clk),
    .D(net274),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _2702_ (.CLK(clknet_leaf_7_clk),
    .D(net74),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_2 _2703_ (.CLK(clknet_leaf_11_clk),
    .D(net267),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfrtp_1 _2704_ (.CLK(clknet_leaf_13_clk),
    .D(net206),
    .RESET_B(net172),
    .Q(\gray_sobel0.gray_scale0.nreset_i ));
 sky130_fd_sc_hd__dfrtp_1 _2705_ (.CLK(clknet_leaf_13_clk),
    .D(net137),
    .RESET_B(net172),
    .Q(\nreset_sync0.r_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2706_ (.CLK(clknet_leaf_11_clk),
    .D(net212),
    .RESET_B(net107),
    .Q(\gray_sobel0.select_sobel_mux ));
 sky130_fd_sc_hd__dfrtp_1 _2707_ (.CLK(clknet_leaf_12_clk),
    .D(net181),
    .RESET_B(net111),
    .Q(\sgnl_sync0.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2708_ (.CLK(clknet_leaf_11_clk),
    .D(net208),
    .RESET_B(net108),
    .Q(\sgnl_sync1.signal_o ));
 sky130_fd_sc_hd__dfrtp_1 _2709_ (.CLK(clknet_leaf_11_clk),
    .D(net189),
    .RESET_B(net108),
    .Q(\sgnl_sync1.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2710_ (.CLK(clknet_leaf_11_clk),
    .D(net216),
    .RESET_B(net108),
    .Q(LFSR_enable_i_sync));
 sky130_fd_sc_hd__dfrtp_1 _2711_ (.CLK(clknet_leaf_11_clk),
    .D(net175),
    .RESET_B(net107),
    .Q(\sgnl_sync2.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2712_ (.CLK(clknet_leaf_11_clk),
    .D(net207),
    .RESET_B(net109),
    .Q(\lfsr0.config_i ));
 sky130_fd_sc_hd__dfrtp_1 _2713_ (.CLK(clknet_leaf_11_clk),
    .D(net183),
    .RESET_B(net108),
    .Q(\sgnl_sync3.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2714_ (.CLK(clknet_leaf_10_clk),
    .D(net213),
    .RESET_B(net108),
    .Q(\lfsr0.lfsr_en_i ));
 sky130_fd_sc_hd__dfrtp_1 _2715_ (.CLK(clknet_leaf_10_clk),
    .D(net191),
    .RESET_B(net108),
    .Q(\sgnl_sync4.signal_sync ));
 sky130_fd_sc_hd__dfrtp_2 _2716_ (.CLK(clknet_leaf_11_clk),
    .D(net214),
    .RESET_B(net108),
    .Q(\sa0.en_i ));
 sky130_fd_sc_hd__dfrtp_1 _2717_ (.CLK(clknet_leaf_12_clk),
    .D(net179),
    .RESET_B(net111),
    .Q(\sgnl_sync5.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2718_ (.CLK(clknet_leaf_11_clk),
    .D(net210),
    .RESET_B(net109),
    .Q(frame_done_i_sync));
 sky130_fd_sc_hd__dfrtp_1 _2719_ (.CLK(clknet_leaf_11_clk),
    .D(net185),
    .RESET_B(net107),
    .Q(\sgnl_sync6.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2720_ (.CLK(clknet_leaf_11_clk),
    .D(net215),
    .RESET_B(net108),
    .Q(lfsr_mode_sel_i_sync));
 sky130_fd_sc_hd__dfrtp_1 _2721_ (.CLK(clknet_leaf_11_clk),
    .D(net177),
    .RESET_B(net107),
    .Q(\sgnl_sync7.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2722_ (.CLK(clknet_leaf_10_clk),
    .D(net209),
    .RESET_B(net108),
    .Q(\sa0.clear_i ));
 sky130_fd_sc_hd__dfrtp_1 _2723_ (.CLK(clknet_leaf_10_clk),
    .D(net187),
    .RESET_B(net108),
    .Q(\sgnl_sync8.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2724_ (.CLK(net141),
    .D(_0002_),
    .RESET_B(_0041_),
    .Q(\spi0.spi0.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2725_ (.CLK(net142),
    .D(_0003_),
    .RESET_B(_0043_),
    .Q(\spi0.spi0.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2726_ (.CLK(net143),
    .D(_0004_),
    .RESET_B(_0045_),
    .Q(\spi0.spi0.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2727_ (.CLK(net144),
    .D(_0005_),
    .RESET_B(_0047_),
    .Q(\spi0.spi0.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2728_ (.CLK(net145),
    .D(_0006_),
    .RESET_B(_0049_),
    .Q(\spi0.spi0.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2729_ (.CLK(net146),
    .D(_0007_),
    .RESET_B(_0051_),
    .Q(\spi0.spi0.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2730_ (.CLK(clknet_2_2__leaf_ui_in[1]),
    .D(net50),
    .RESET_B(_0053_),
    .Q(\spi0.signal_sync1.async_signal_i ));
 sky130_fd_sc_hd__dfrtp_1 _2731_ (.CLK(net147),
    .D(_0009_),
    .RESET_B(_0054_),
    .Q(\spi0.spi0.sdo_register[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2732_ (.CLK(net148),
    .D(_0020_),
    .RESET_B(_0056_),
    .Q(\spi0.spi0.sdo_register[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2733_ (.CLK(net149),
    .D(_0025_),
    .RESET_B(_0058_),
    .Q(\spi0.spi0.sdo_register[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2734_ (.CLK(net150),
    .D(_0026_),
    .RESET_B(_0060_),
    .Q(\spi0.spi0.sdo_register[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2735_ (.CLK(net151),
    .D(_0027_),
    .RESET_B(_0062_),
    .Q(\spi0.spi0.sdo_register[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2736_ (.CLK(net152),
    .D(_0028_),
    .RESET_B(_0064_),
    .Q(\spi0.spi0.sdo_register[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2737_ (.CLK(net153),
    .D(_0029_),
    .RESET_B(_0066_),
    .Q(\spi0.spi0.sdo_register[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2738_ (.CLK(net154),
    .D(_0030_),
    .RESET_B(_0068_),
    .Q(\spi0.spi0.sdo_register[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2739_ (.CLK(net155),
    .D(_0031_),
    .RESET_B(_0070_),
    .Q(\spi0.spi0.sdo_register[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2740_ (.CLK(net156),
    .D(_0032_),
    .RESET_B(_0072_),
    .Q(\spi0.spi0.sdo_register[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2741_ (.CLK(net157),
    .D(_0010_),
    .RESET_B(_0074_),
    .Q(\spi0.spi0.sdo_register[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2742_ (.CLK(net158),
    .D(_0011_),
    .RESET_B(_0076_),
    .Q(\spi0.spi0.sdo_register[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2743_ (.CLK(net159),
    .D(_0012_),
    .RESET_B(_0078_),
    .Q(\spi0.spi0.sdo_register[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2744_ (.CLK(net160),
    .D(_0013_),
    .RESET_B(_0080_),
    .Q(\spi0.spi0.sdo_register[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2745_ (.CLK(net161),
    .D(_0014_),
    .RESET_B(_0082_),
    .Q(\spi0.spi0.sdo_register[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2746_ (.CLK(net162),
    .D(_0015_),
    .RESET_B(_0084_),
    .Q(\spi0.spi0.sdo_register[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2747_ (.CLK(net163),
    .D(_0016_),
    .RESET_B(_0086_),
    .Q(\spi0.spi0.sdo_register[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2748_ (.CLK(net164),
    .D(_0017_),
    .RESET_B(_0088_),
    .Q(\spi0.spi0.sdo_register[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2749_ (.CLK(net165),
    .D(_0018_),
    .RESET_B(_0090_),
    .Q(\spi0.spi0.sdo_register[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2750_ (.CLK(net166),
    .D(_0019_),
    .RESET_B(_0092_),
    .Q(\spi0.spi0.sdo_register[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2751_ (.CLK(net167),
    .D(_0021_),
    .RESET_B(_0094_),
    .Q(\spi0.spi0.sdo_register[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2752_ (.CLK(net168),
    .D(_0022_),
    .RESET_B(_0096_),
    .Q(\spi0.spi0.sdo_register[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2753_ (.CLK(net169),
    .D(_0023_),
    .RESET_B(_0098_),
    .Q(\spi0.spi0.sdo_register[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2754_ (.CLK(net170),
    .D(_0024_),
    .RESET_B(_0100_),
    .Q(\spi0.spi0.sdo_o ));
 sky130_fd_sc_hd__dfrtp_1 _2755_ (.CLK(clknet_leaf_20_clk),
    .D(_0126_),
    .RESET_B(net79),
    .Q(\input_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2756_ (.CLK(clknet_leaf_20_clk),
    .D(_0127_),
    .RESET_B(net78),
    .Q(\input_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2757_ (.CLK(clknet_leaf_20_clk),
    .D(_0128_),
    .RESET_B(net79),
    .Q(\input_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2758_ (.CLK(clknet_leaf_19_clk),
    .D(_0129_),
    .RESET_B(net84),
    .Q(\input_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2759_ (.CLK(clknet_leaf_19_clk),
    .D(_0130_),
    .RESET_B(net85),
    .Q(\input_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2760_ (.CLK(clknet_leaf_2_clk),
    .D(_0131_),
    .RESET_B(net98),
    .Q(\input_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2761_ (.CLK(clknet_leaf_9_clk),
    .D(_0132_),
    .RESET_B(net98),
    .Q(\input_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2762_ (.CLK(clknet_leaf_9_clk),
    .D(_0133_),
    .RESET_B(net98),
    .Q(\input_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2763_ (.CLK(clknet_leaf_4_clk),
    .D(_0134_),
    .RESET_B(net93),
    .Q(\input_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2764_ (.CLK(clknet_leaf_0_clk),
    .D(_0135_),
    .RESET_B(net82),
    .Q(\input_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2765_ (.CLK(clknet_leaf_23_clk),
    .D(_0136_),
    .RESET_B(net81),
    .Q(\input_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2766_ (.CLK(clknet_leaf_23_clk),
    .D(_0137_),
    .RESET_B(net81),
    .Q(\input_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2767_ (.CLK(clknet_leaf_23_clk),
    .D(_0138_),
    .RESET_B(net80),
    .Q(\input_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2768_ (.CLK(clknet_leaf_23_clk),
    .D(_0139_),
    .RESET_B(net80),
    .Q(\input_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2769_ (.CLK(clknet_leaf_23_clk),
    .D(_0140_),
    .RESET_B(net80),
    .Q(\input_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2770_ (.CLK(clknet_leaf_23_clk),
    .D(_0141_),
    .RESET_B(net80),
    .Q(\input_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2771_ (.CLK(clknet_leaf_8_clk),
    .D(_0142_),
    .RESET_B(net97),
    .Q(\input_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2772_ (.CLK(clknet_leaf_4_clk),
    .D(_0143_),
    .RESET_B(net94),
    .Q(\input_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2773_ (.CLK(clknet_leaf_4_clk),
    .D(_0144_),
    .RESET_B(net94),
    .Q(\input_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2774_ (.CLK(clknet_leaf_4_clk),
    .D(_0145_),
    .RESET_B(net93),
    .Q(\input_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2775_ (.CLK(clknet_leaf_4_clk),
    .D(_0146_),
    .RESET_B(net93),
    .Q(\input_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2776_ (.CLK(clknet_leaf_0_clk),
    .D(_0147_),
    .RESET_B(net82),
    .Q(\input_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2777_ (.CLK(clknet_leaf_23_clk),
    .D(_0148_),
    .RESET_B(net81),
    .Q(\input_data[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2778_ (.CLK(clknet_leaf_0_clk),
    .D(_0149_),
    .RESET_B(net82),
    .Q(\input_data[23] ));
 sky130_fd_sc_hd__dfrtp_2 _2779_ (.CLK(clknet_2_3__leaf_ui_in[1]),
    .D(net195),
    .RESET_B(_0102_),
    .Q(\spi0.spi0.data_rx_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2780_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net279),
    .RESET_B(_0103_),
    .Q(\spi0.spi0.data_rx_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2781_ (.CLK(clknet_2_2__leaf_ui_in[1]),
    .D(net211),
    .RESET_B(_0104_),
    .Q(\spi0.spi0.data_rx_o[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2782_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net242),
    .RESET_B(_0105_),
    .Q(\spi0.spi0.data_rx_o[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2783_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net228),
    .RESET_B(_0106_),
    .Q(\spi0.spi0.data_rx_o[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2784_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net230),
    .RESET_B(_0107_),
    .Q(\spi0.spi0.data_rx_o[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2785_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net236),
    .RESET_B(_0108_),
    .Q(\spi0.spi0.data_rx_o[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2786_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net218),
    .RESET_B(_0109_),
    .Q(\spi0.spi0.data_rx_o[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2787_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net223),
    .RESET_B(_0110_),
    .Q(\spi0.spi0.data_rx_o[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2788_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net232),
    .RESET_B(_0111_),
    .Q(\spi0.spi0.data_rx_o[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2789_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net235),
    .RESET_B(_0112_),
    .Q(\spi0.spi0.data_rx_o[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2790_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net229),
    .RESET_B(_0113_),
    .Q(\spi0.spi0.data_rx_o[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2791_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net233),
    .RESET_B(_0114_),
    .Q(\spi0.spi0.data_rx_o[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2792_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net226),
    .RESET_B(_0115_),
    .Q(\spi0.spi0.data_rx_o[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2793_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net221),
    .RESET_B(_0116_),
    .Q(\spi0.spi0.data_rx_o[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2794_ (.CLK(clknet_2_0__leaf_ui_in[1]),
    .D(net220),
    .RESET_B(_0117_),
    .Q(\spi0.spi0.data_rx_o[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2795_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net231),
    .RESET_B(_0118_),
    .Q(\spi0.spi0.data_rx_o[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2796_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net227),
    .RESET_B(_0119_),
    .Q(\spi0.spi0.data_rx_o[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2797_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net225),
    .RESET_B(_0120_),
    .Q(\spi0.spi0.data_rx_o[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2798_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net219),
    .RESET_B(_0121_),
    .Q(\spi0.spi0.data_rx_o[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2799_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net238),
    .RESET_B(_0122_),
    .Q(\spi0.spi0.data_rx_o[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2800_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net239),
    .RESET_B(_0123_),
    .Q(\spi0.spi0.data_rx_o[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2801_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net217),
    .RESET_B(_0124_),
    .Q(\spi0.spi0.data_rx_o[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2802_ (.CLK(clknet_2_1__leaf_ui_in[1]),
    .D(net224),
    .RESET_B(_0125_),
    .Q(\spi0.spi0.data_rx_o[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2803_ (.CLK(clknet_leaf_4_clk),
    .D(\spi0.signal_sync1.async_signal_i ),
    .RESET_B(net94),
    .Q(\spi0.signal_sync1.signal_sync ));
 sky130_fd_sc_hd__dfrtp_1 _2804_ (.CLK(clknet_leaf_4_clk),
    .D(net205),
    .RESET_B(net94),
    .Q(\spi0.rxtx_done ));
 sky130_fd_sc_hd__dfrtp_1 _2805_ (.CLK(clknet_leaf_8_clk),
    .D(net64),
    .RESET_B(net99),
    .Q(in_data_rdy));
 sky130_fd_sc_hd__dfrtp_1 _2806_ (.CLK(clknet_leaf_8_clk),
    .D(_0150_),
    .RESET_B(net102),
    .Q(\spi0.data_tx[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2807_ (.CLK(clknet_leaf_8_clk),
    .D(_0151_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2808_ (.CLK(clknet_leaf_8_clk),
    .D(_0152_),
    .RESET_B(net102),
    .Q(\spi0.data_tx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2809_ (.CLK(clknet_leaf_7_clk),
    .D(_0153_),
    .RESET_B(net102),
    .Q(\spi0.data_tx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2810_ (.CLK(clknet_leaf_11_clk),
    .D(_0154_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2811_ (.CLK(clknet_leaf_7_clk),
    .D(_0155_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2812_ (.CLK(clknet_leaf_7_clk),
    .D(_0156_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2813_ (.CLK(clknet_leaf_7_clk),
    .D(_0157_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2814_ (.CLK(clknet_leaf_6_clk),
    .D(_0158_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2815_ (.CLK(clknet_leaf_6_clk),
    .D(_0159_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2816_ (.CLK(clknet_leaf_7_clk),
    .D(_0160_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2817_ (.CLK(clknet_leaf_7_clk),
    .D(_0161_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2818_ (.CLK(clknet_leaf_7_clk),
    .D(_0162_),
    .RESET_B(net103),
    .Q(\spi0.data_tx[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2819_ (.CLK(clknet_leaf_6_clk),
    .D(_0163_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2820_ (.CLK(clknet_leaf_6_clk),
    .D(_0164_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2821_ (.CLK(clknet_leaf_6_clk),
    .D(_0165_),
    .RESET_B(net102),
    .Q(\spi0.data_tx[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2822_ (.CLK(clknet_leaf_6_clk),
    .D(_0166_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2823_ (.CLK(clknet_leaf_5_clk),
    .D(_0167_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2824_ (.CLK(clknet_leaf_4_clk),
    .D(_0168_),
    .RESET_B(net100),
    .Q(\spi0.data_tx[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2825_ (.CLK(clknet_leaf_5_clk),
    .D(_0169_),
    .RESET_B(net100),
    .Q(\spi0.data_tx[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2826_ (.CLK(clknet_leaf_4_clk),
    .D(_0170_),
    .RESET_B(net100),
    .Q(\spi0.data_tx[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2827_ (.CLK(clknet_leaf_5_clk),
    .D(_0171_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2828_ (.CLK(clknet_leaf_6_clk),
    .D(_0172_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2829_ (.CLK(clknet_leaf_6_clk),
    .D(_0173_),
    .RESET_B(net101),
    .Q(\spi0.data_tx[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2830_ (.CLK(clknet_leaf_8_clk),
    .D(_0174_),
    .RESET_B(net99),
    .Q(\sa0.signature_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2831_ (.CLK(clknet_leaf_8_clk),
    .D(_0175_),
    .RESET_B(net97),
    .Q(\sa0.signature_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2832_ (.CLK(clknet_leaf_8_clk),
    .D(_0176_),
    .RESET_B(net97),
    .Q(\sa0.signature_o[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2833_ (.CLK(clknet_leaf_9_clk),
    .D(_0177_),
    .RESET_B(net105),
    .Q(\sa0.signature_o[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2834_ (.CLK(clknet_leaf_9_clk),
    .D(_0178_),
    .RESET_B(net105),
    .Q(\sa0.signature_o[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2835_ (.CLK(clknet_leaf_8_clk),
    .D(_0179_),
    .RESET_B(net99),
    .Q(\sa0.signature_o[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2836_ (.CLK(clknet_leaf_8_clk),
    .D(_0180_),
    .RESET_B(net102),
    .Q(\sa0.signature_o[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2837_ (.CLK(clknet_leaf_8_clk),
    .D(_0181_),
    .RESET_B(net97),
    .Q(\sa0.signature_o[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2838_ (.CLK(clknet_leaf_3_clk),
    .D(_0182_),
    .RESET_B(net97),
    .Q(\sa0.signature_o[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2839_ (.CLK(clknet_leaf_3_clk),
    .D(_0183_),
    .RESET_B(net97),
    .Q(\sa0.signature_o[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2840_ (.CLK(clknet_leaf_3_clk),
    .D(_0184_),
    .RESET_B(net102),
    .Q(\sa0.signature_o[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2841_ (.CLK(clknet_leaf_8_clk),
    .D(_0185_),
    .RESET_B(net102),
    .Q(\sa0.signature_o[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2842_ (.CLK(clknet_leaf_8_clk),
    .D(net371),
    .RESET_B(net102),
    .Q(\sa0.signature_o[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2843_ (.CLK(clknet_leaf_8_clk),
    .D(net401),
    .RESET_B(net102),
    .Q(\sa0.signature_o[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2844_ (.CLK(clknet_leaf_6_clk),
    .D(_0188_),
    .RESET_B(net100),
    .Q(\sa0.signature_o[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2845_ (.CLK(clknet_leaf_6_clk),
    .D(net378),
    .RESET_B(net100),
    .Q(\sa0.signature_o[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2846_ (.CLK(clknet_leaf_5_clk),
    .D(net381),
    .RESET_B(net100),
    .Q(\sa0.signature_o[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2847_ (.CLK(clknet_leaf_6_clk),
    .D(_0191_),
    .RESET_B(net100),
    .Q(\sa0.signature_o[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2848_ (.CLK(clknet_leaf_5_clk),
    .D(net361),
    .RESET_B(net100),
    .Q(\sa0.signature_o[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2849_ (.CLK(clknet_leaf_5_clk),
    .D(net383),
    .RESET_B(net100),
    .Q(\sa0.signature_o[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2850_ (.CLK(clknet_leaf_5_clk),
    .D(net387),
    .RESET_B(net100),
    .Q(\sa0.signature_o[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2851_ (.CLK(clknet_leaf_4_clk),
    .D(_0195_),
    .RESET_B(net94),
    .Q(\sa0.signature_o[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2852_ (.CLK(clknet_leaf_4_clk),
    .D(net389),
    .RESET_B(net94),
    .Q(\sa0.signature_o[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2853_ (.CLK(clknet_leaf_5_clk),
    .D(net318),
    .RESET_B(net95),
    .Q(\sa0.signature_o[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2854_ (.CLK(clknet_leaf_4_clk),
    .D(net222),
    .RESET_B(net94),
    .Q(\spi0.rxtx_done_reg ));
 sky130_fd_sc_hd__dfrtp_1 _2855_ (.CLK(clknet_leaf_12_clk),
    .D(\gray_sobel0.sobel0.next[0] ),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.fsm_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2856_ (.CLK(clknet_leaf_12_clk),
    .D(net47),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.fsm_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2857_ (.CLK(clknet_leaf_9_clk),
    .D(net373),
    .RESET_B(net109),
    .Q(\gray_sobel0.px_rdy_o_sobel ));
 sky130_fd_sc_hd__dfrtp_1 _2858_ (.CLK(clknet_leaf_16_clk),
    .D(_0198_),
    .RESET_B(net88),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2859_ (.CLK(clknet_leaf_16_clk),
    .D(_0199_),
    .RESET_B(net88),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2860_ (.CLK(clknet_leaf_16_clk),
    .D(_0200_),
    .RESET_B(net88),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2861_ (.CLK(clknet_leaf_18_clk),
    .D(_0201_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2862_ (.CLK(clknet_leaf_15_clk),
    .D(_0202_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2863_ (.CLK(clknet_leaf_15_clk),
    .D(_0203_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2864_ (.CLK(clknet_leaf_14_clk),
    .D(_0204_),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2865_ (.CLK(clknet_leaf_10_clk),
    .D(_0205_),
    .RESET_B(net109),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2866_ (.CLK(clknet_leaf_9_clk),
    .D(_0206_),
    .RESET_B(net104),
    .Q(\gray_sobel0.out_px_sobel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2867_ (.CLK(clknet_leaf_15_clk),
    .D(_0207_),
    .RESET_B(net104),
    .Q(\gray_sobel0.out_px_sobel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2868_ (.CLK(clknet_leaf_15_clk),
    .D(_0208_),
    .RESET_B(net104),
    .Q(\gray_sobel0.out_px_sobel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2869_ (.CLK(clknet_leaf_9_clk),
    .D(_0209_),
    .RESET_B(net104),
    .Q(\gray_sobel0.out_px_sobel[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2870_ (.CLK(clknet_leaf_15_clk),
    .D(_0210_),
    .RESET_B(net104),
    .Q(\gray_sobel0.out_px_sobel[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2871_ (.CLK(clknet_leaf_15_clk),
    .D(_0211_),
    .RESET_B(net98),
    .Q(\gray_sobel0.out_px_sobel[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2872_ (.CLK(clknet_leaf_15_clk),
    .D(_0212_),
    .RESET_B(net104),
    .Q(\gray_sobel0.out_px_sobel[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2873_ (.CLK(clknet_leaf_15_clk),
    .D(_0213_),
    .RESET_B(net104),
    .Q(\gray_sobel0.out_px_sobel[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2874_ (.CLK(clknet_leaf_21_clk),
    .D(_0214_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2875_ (.CLK(clknet_leaf_21_clk),
    .D(_0215_),
    .RESET_B(net78),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2876_ (.CLK(clknet_leaf_17_clk),
    .D(_0216_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2877_ (.CLK(clknet_leaf_18_clk),
    .D(_0217_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2878_ (.CLK(clknet_leaf_18_clk),
    .D(_0218_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2879_ (.CLK(clknet_leaf_19_clk),
    .D(_0219_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2880_ (.CLK(clknet_leaf_9_clk),
    .D(_0220_),
    .RESET_B(net104),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2881_ (.CLK(clknet_leaf_9_clk),
    .D(_0221_),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2882_ (.CLK(clknet_leaf_12_clk),
    .D(_0222_),
    .RESET_B(net109),
    .Q(\gray_sobel0.sobel0.counter_sobel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2883_ (.CLK(clknet_leaf_10_clk),
    .D(_0223_),
    .RESET_B(net109),
    .Q(\gray_sobel0.sobel0.counter_sobel[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2884_ (.CLK(clknet_leaf_10_clk),
    .D(_0224_),
    .RESET_B(net107),
    .Q(\gray_sobel0.sobel0.counter_sobel[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2885_ (.CLK(clknet_leaf_11_clk),
    .D(_0225_),
    .RESET_B(net107),
    .Q(\gray_sobel0.sobel0.counter_sobel[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2886_ (.CLK(clknet_leaf_9_clk),
    .D(net28),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.px_ready ));
 sky130_fd_sc_hd__dfrtp_1 _2887_ (.CLK(clknet_leaf_16_clk),
    .D(_0226_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2888_ (.CLK(clknet_leaf_17_clk),
    .D(_0227_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2889_ (.CLK(clknet_leaf_17_clk),
    .D(_0228_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2890_ (.CLK(clknet_leaf_18_clk),
    .D(_0229_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2891_ (.CLK(clknet_leaf_18_clk),
    .D(_0230_),
    .RESET_B(net91),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2892_ (.CLK(clknet_leaf_15_clk),
    .D(_0231_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2893_ (.CLK(clknet_leaf_15_clk),
    .D(_0232_),
    .RESET_B(net104),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[6] ));
 sky130_fd_sc_hd__dfrtp_2 _2894_ (.CLK(clknet_leaf_10_clk),
    .D(_0233_),
    .RESET_B(net106),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i6[7] ));
 sky130_fd_sc_hd__dfrtp_2 _2895_ (.CLK(clknet_leaf_11_clk),
    .D(_0234_),
    .RESET_B(net107),
    .Q(\gray_sobel0.sobel0.counter_pixels[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2896_ (.CLK(clknet_leaf_11_clk),
    .D(_0235_),
    .RESET_B(net107),
    .Q(\gray_sobel0.sobel0.counter_pixels[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2897_ (.CLK(clknet_leaf_11_clk),
    .D(_0236_),
    .RESET_B(net107),
    .Q(\gray_sobel0.sobel0.counter_pixels[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2898_ (.CLK(clknet_leaf_11_clk),
    .D(_0237_),
    .RESET_B(net107),
    .Q(\gray_sobel0.sobel0.counter_pixels[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2899_ (.CLK(clknet_leaf_12_clk),
    .D(_0238_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2900_ (.CLK(clknet_leaf_11_clk),
    .D(_0239_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2901_ (.CLK(clknet_leaf_12_clk),
    .D(_0240_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2902_ (.CLK(clknet_leaf_12_clk),
    .D(_0241_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2903_ (.CLK(clknet_leaf_13_clk),
    .D(_0242_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2904_ (.CLK(clknet_leaf_13_clk),
    .D(_0243_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2905_ (.CLK(clknet_leaf_13_clk),
    .D(_0244_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2906_ (.CLK(clknet_leaf_13_clk),
    .D(_0245_),
    .RESET_B(net112),
    .Q(\gray_sobel0.sobel0.counter_pixels[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2907_ (.CLK(clknet_leaf_13_clk),
    .D(_0246_),
    .RESET_B(net112),
    .Q(\gray_sobel0.sobel0.counter_pixels[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2908_ (.CLK(clknet_leaf_13_clk),
    .D(_0247_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.counter_pixels[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2909_ (.CLK(clknet_leaf_13_clk),
    .D(_0248_),
    .RESET_B(net112),
    .Q(\gray_sobel0.sobel0.counter_pixels[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2910_ (.CLK(clknet_leaf_13_clk),
    .D(_0249_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.counter_pixels[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2911_ (.CLK(clknet_leaf_12_clk),
    .D(_0250_),
    .RESET_B(net111),
    .Q(\gray_sobel0.sobel0.counter_pixels[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2912_ (.CLK(clknet_leaf_12_clk),
    .D(_0251_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.counter_pixels[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2913_ (.CLK(clknet_leaf_12_clk),
    .D(_0252_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.counter_pixels[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2914_ (.CLK(clknet_leaf_14_clk),
    .D(_0253_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.counter_pixels[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2915_ (.CLK(clknet_leaf_13_clk),
    .D(_0254_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.counter_pixels[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2916_ (.CLK(clknet_leaf_13_clk),
    .D(_0255_),
    .RESET_B(net112),
    .Q(\gray_sobel0.sobel0.counter_pixels[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2917_ (.CLK(clknet_leaf_13_clk),
    .D(_0256_),
    .RESET_B(net112),
    .Q(\gray_sobel0.sobel0.counter_pixels[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2918_ (.CLK(clknet_leaf_13_clk),
    .D(_0257_),
    .RESET_B(net112),
    .Q(\gray_sobel0.sobel0.counter_pixels[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2919_ (.CLK(clknet_leaf_16_clk),
    .D(_0258_),
    .RESET_B(net91),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2920_ (.CLK(clknet_leaf_16_clk),
    .D(_0259_),
    .RESET_B(net91),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2921_ (.CLK(clknet_leaf_16_clk),
    .D(_0260_),
    .RESET_B(net88),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2922_ (.CLK(clknet_leaf_18_clk),
    .D(_0261_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2923_ (.CLK(clknet_leaf_15_clk),
    .D(_0262_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2924_ (.CLK(clknet_leaf_15_clk),
    .D(_0263_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2925_ (.CLK(clknet_leaf_14_clk),
    .D(_0264_),
    .RESET_B(net113),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2926_ (.CLK(clknet_leaf_12_clk),
    .D(_0265_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2927_ (.CLK(clknet_leaf_17_clk),
    .D(_0266_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2928_ (.CLK(clknet_leaf_21_clk),
    .D(_0267_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2929_ (.CLK(clknet_leaf_17_clk),
    .D(_0268_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2930_ (.CLK(clknet_leaf_18_clk),
    .D(_0269_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2931_ (.CLK(clknet_leaf_18_clk),
    .D(_0270_),
    .RESET_B(net91),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2932_ (.CLK(clknet_leaf_19_clk),
    .D(_0271_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2933_ (.CLK(clknet_leaf_9_clk),
    .D(_0272_),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2934_ (.CLK(clknet_leaf_9_clk),
    .D(_0273_),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2935_ (.CLK(clknet_leaf_16_clk),
    .D(_0274_),
    .RESET_B(net88),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2936_ (.CLK(clknet_leaf_16_clk),
    .D(_0275_),
    .RESET_B(net88),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2937_ (.CLK(clknet_leaf_17_clk),
    .D(_0276_),
    .RESET_B(net88),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2938_ (.CLK(clknet_leaf_18_clk),
    .D(_0277_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2939_ (.CLK(clknet_leaf_18_clk),
    .D(_0278_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2940_ (.CLK(clknet_leaf_15_clk),
    .D(_0279_),
    .RESET_B(net106),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2941_ (.CLK(clknet_leaf_14_clk),
    .D(_0280_),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2942_ (.CLK(clknet_leaf_10_clk),
    .D(_0281_),
    .RESET_B(net109),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2943_ (.CLK(clknet_leaf_16_clk),
    .D(_0282_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2944_ (.CLK(clknet_leaf_16_clk),
    .D(_0283_),
    .RESET_B(net91),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2945_ (.CLK(clknet_leaf_18_clk),
    .D(_0284_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2946_ (.CLK(clknet_leaf_18_clk),
    .D(_0285_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2947_ (.CLK(clknet_leaf_15_clk),
    .D(_0286_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2948_ (.CLK(clknet_leaf_15_clk),
    .D(_0287_),
    .RESET_B(net106),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[5] ));
 sky130_fd_sc_hd__dfrtp_4 _2949_ (.CLK(clknet_leaf_14_clk),
    .D(_0288_),
    .RESET_B(net113),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2950_ (.CLK(clknet_leaf_12_clk),
    .D(_0289_),
    .RESET_B(net110),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2951_ (.CLK(clknet_leaf_17_clk),
    .D(_0290_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2952_ (.CLK(clknet_leaf_17_clk),
    .D(_0291_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2953_ (.CLK(clknet_leaf_20_clk),
    .D(_0292_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2954_ (.CLK(clknet_leaf_18_clk),
    .D(_0293_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2955_ (.CLK(clknet_leaf_18_clk),
    .D(_0294_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2956_ (.CLK(clknet_leaf_19_clk),
    .D(_0295_),
    .RESET_B(net90),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2957_ (.CLK(clknet_leaf_9_clk),
    .D(_0296_),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2958_ (.CLK(clknet_leaf_9_clk),
    .D(_0297_),
    .RESET_B(net105),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2959_ (.CLK(clknet_leaf_20_clk),
    .D(_0033_),
    .RESET_B(net79),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2960_ (.CLK(clknet_leaf_20_clk),
    .D(_0034_),
    .RESET_B(net78),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2961_ (.CLK(clknet_leaf_21_clk),
    .D(_0035_),
    .RESET_B(net78),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2962_ (.CLK(clknet_leaf_21_clk),
    .D(_0036_),
    .RESET_B(net78),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2963_ (.CLK(clknet_leaf_21_clk),
    .D(_0037_),
    .RESET_B(net78),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2964_ (.CLK(clknet_leaf_21_clk),
    .D(_0038_),
    .RESET_B(net78),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2965_ (.CLK(clknet_leaf_22_clk),
    .D(_0039_),
    .RESET_B(net78),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2966_ (.CLK(clknet_leaf_22_clk),
    .D(_0040_),
    .RESET_B(net78),
    .Q(\gray_sobel0.gray_scale0.out_px_gray_o[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2967_ (.CLK(clknet_leaf_10_clk),
    .D(\gray_sobel0.gray_scale0.px_rdy_i ),
    .RESET_B(net109),
    .Q(\gray_sobel0.gray_scale0.px_rdy_o ));
 sky130_fd_sc_hd__dfrtp_1 _2968_ (.CLK(clknet_leaf_8_clk),
    .D(in_lfsr_rdy),
    .RESET_B(net102),
    .Q(\lfsr0.config_done_o ));
 sky130_fd_sc_hd__dfrtp_1 _2969_ (.CLK(clknet_leaf_10_clk),
    .D(_0000_),
    .RESET_B(net109),
    .Q(\lfsr0.lfsr_rdy_o ));
 sky130_fd_sc_hd__dfrtp_2 _2970_ (.CLK(clknet_leaf_1_clk),
    .D(_0298_),
    .RESET_B(net84),
    .Q(\lfsr0.lfsr_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2971_ (.CLK(clknet_leaf_20_clk),
    .D(_0299_),
    .RESET_B(net84),
    .Q(\lfsr0.lfsr_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2972_ (.CLK(clknet_leaf_19_clk),
    .D(_0300_),
    .RESET_B(net84),
    .Q(\lfsr0.lfsr_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _2973_ (.CLK(clknet_leaf_19_clk),
    .D(_0301_),
    .RESET_B(net84),
    .Q(\lfsr0.lfsr_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _2974_ (.CLK(clknet_leaf_19_clk),
    .D(_0302_),
    .RESET_B(net85),
    .Q(\lfsr0.lfsr_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2975_ (.CLK(clknet_leaf_1_clk),
    .D(_0303_),
    .RESET_B(net85),
    .Q(\lfsr0.lfsr_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _2976_ (.CLK(clknet_leaf_2_clk),
    .D(_0304_),
    .RESET_B(net98),
    .Q(\lfsr0.lfsr_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2977_ (.CLK(clknet_leaf_3_clk),
    .D(_0305_),
    .RESET_B(net98),
    .Q(\lfsr0.lfsr_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2978_ (.CLK(clknet_leaf_3_clk),
    .D(_0306_),
    .RESET_B(net98),
    .Q(\lfsr0.lfsr_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2979_ (.CLK(clknet_leaf_0_clk),
    .D(_0307_),
    .RESET_B(net83),
    .Q(\lfsr0.lfsr_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2980_ (.CLK(clknet_leaf_1_clk),
    .D(_0308_),
    .RESET_B(net81),
    .Q(\lfsr0.lfsr_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _2981_ (.CLK(clknet_leaf_1_clk),
    .D(_0309_),
    .RESET_B(net84),
    .Q(\lfsr0.lfsr_out[11] ));
 sky130_fd_sc_hd__dfrtp_2 _2982_ (.CLK(clknet_leaf_20_clk),
    .D(_0310_),
    .RESET_B(net79),
    .Q(\lfsr0.lfsr_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _2983_ (.CLK(clknet_leaf_23_clk),
    .D(_0311_),
    .RESET_B(net81),
    .Q(\lfsr0.lfsr_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2984_ (.CLK(clknet_leaf_23_clk),
    .D(_0312_),
    .RESET_B(net83),
    .Q(\lfsr0.lfsr_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2985_ (.CLK(clknet_leaf_0_clk),
    .D(_0313_),
    .RESET_B(net82),
    .Q(\lfsr0.lfsr_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _2986_ (.CLK(clknet_leaf_3_clk),
    .D(_0314_),
    .RESET_B(net95),
    .Q(\lfsr0.lfsr_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2987_ (.CLK(clknet_leaf_3_clk),
    .D(_0315_),
    .RESET_B(net95),
    .Q(\lfsr0.lfsr_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2988_ (.CLK(clknet_leaf_3_clk),
    .D(_0316_),
    .RESET_B(net95),
    .Q(\lfsr0.lfsr_out[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2989_ (.CLK(clknet_leaf_4_clk),
    .D(_0317_),
    .RESET_B(net93),
    .Q(\lfsr0.lfsr_out[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2990_ (.CLK(clknet_leaf_0_clk),
    .D(_0318_),
    .RESET_B(net93),
    .Q(\lfsr0.lfsr_out[20] ));
 sky130_fd_sc_hd__dfrtp_1 _2991_ (.CLK(clknet_leaf_0_clk),
    .D(_0319_),
    .RESET_B(net83),
    .Q(\lfsr0.lfsr_out[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2992_ (.CLK(clknet_leaf_23_clk),
    .D(_0320_),
    .RESET_B(net81),
    .Q(\lfsr0.lfsr_out[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2993_ (.CLK(clknet_leaf_0_clk),
    .D(_0321_),
    .RESET_B(net82),
    .Q(\lfsr0.lfsr_out[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2994_ (.CLK(clknet_leaf_16_clk),
    .D(_0322_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2995_ (.CLK(clknet_leaf_16_clk),
    .D(_0323_),
    .RESET_B(net86),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2996_ (.CLK(clknet_leaf_17_clk),
    .D(_0324_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2997_ (.CLK(clknet_leaf_17_clk),
    .D(_0325_),
    .RESET_B(net87),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2998_ (.CLK(clknet_leaf_18_clk),
    .D(_0326_),
    .RESET_B(net89),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2999_ (.CLK(clknet_leaf_15_clk),
    .D(_0327_),
    .RESET_B(net106),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3000_ (.CLK(clknet_leaf_15_clk),
    .D(_0328_),
    .RESET_B(net104),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3001_ (.CLK(clknet_leaf_9_clk),
    .D(_0329_),
    .RESET_B(net106),
    .Q(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3002_ (.CLK(clknet_leaf_1_clk),
    .D(_0330_),
    .RESET_B(net85),
    .Q(\lfsr0.seed_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3003_ (.CLK(clknet_leaf_19_clk),
    .D(net325),
    .RESET_B(net84),
    .Q(\lfsr0.seed_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3004_ (.CLK(clknet_leaf_20_clk),
    .D(net351),
    .RESET_B(net79),
    .Q(\lfsr0.seed_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3005_ (.CLK(clknet_leaf_18_clk),
    .D(net376),
    .RESET_B(net89),
    .Q(\lfsr0.seed_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3006_ (.CLK(clknet_leaf_19_clk),
    .D(net353),
    .RESET_B(net85),
    .Q(\lfsr0.seed_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3007_ (.CLK(clknet_leaf_2_clk),
    .D(net333),
    .RESET_B(net85),
    .Q(\lfsr0.seed_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3008_ (.CLK(clknet_leaf_2_clk),
    .D(net329),
    .RESET_B(net98),
    .Q(\lfsr0.seed_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3009_ (.CLK(clknet_leaf_2_clk),
    .D(_0337_),
    .RESET_B(net97),
    .Q(\lfsr0.seed_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3010_ (.CLK(clknet_leaf_3_clk),
    .D(_0338_),
    .RESET_B(net96),
    .Q(\lfsr0.seed_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3011_ (.CLK(clknet_leaf_3_clk),
    .D(_0339_),
    .RESET_B(net93),
    .Q(\lfsr0.seed_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3012_ (.CLK(clknet_leaf_1_clk),
    .D(_0340_),
    .RESET_B(net83),
    .Q(\lfsr0.seed_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3013_ (.CLK(clknet_leaf_20_clk),
    .D(_0341_),
    .RESET_B(net84),
    .Q(\lfsr0.seed_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _3014_ (.CLK(clknet_leaf_22_clk),
    .D(_0342_),
    .RESET_B(net78),
    .Q(\lfsr0.seed_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _3015_ (.CLK(clknet_leaf_23_clk),
    .D(net337),
    .RESET_B(net80),
    .Q(\lfsr0.seed_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _3016_ (.CLK(clknet_leaf_23_clk),
    .D(net355),
    .RESET_B(net80),
    .Q(\lfsr0.seed_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _3017_ (.CLK(clknet_leaf_0_clk),
    .D(_0345_),
    .RESET_B(net82),
    .Q(\lfsr0.seed_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _3018_ (.CLK(clknet_leaf_3_clk),
    .D(net369),
    .RESET_B(net97),
    .Q(\lfsr0.seed_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _3019_ (.CLK(clknet_leaf_3_clk),
    .D(net342),
    .RESET_B(net94),
    .Q(\lfsr0.seed_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _3020_ (.CLK(clknet_leaf_4_clk),
    .D(net340),
    .RESET_B(net94),
    .Q(\lfsr0.seed_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _3021_ (.CLK(clknet_leaf_4_clk),
    .D(net357),
    .RESET_B(net93),
    .Q(\lfsr0.seed_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _3022_ (.CLK(clknet_leaf_4_clk),
    .D(net323),
    .RESET_B(net93),
    .Q(\lfsr0.seed_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _3023_ (.CLK(clknet_leaf_0_clk),
    .D(net363),
    .RESET_B(net82),
    .Q(\lfsr0.seed_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _3024_ (.CLK(clknet_leaf_23_clk),
    .D(net345),
    .RESET_B(net81),
    .Q(\lfsr0.seed_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _3025_ (.CLK(clknet_leaf_0_clk),
    .D(net347),
    .RESET_B(net82),
    .Q(\lfsr0.seed_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _3026_ (.CLK(clknet_leaf_1_clk),
    .D(_0354_),
    .RESET_B(net85),
    .Q(\lfsr0.stop_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3027_ (.CLK(clknet_leaf_19_clk),
    .D(net398),
    .RESET_B(net84),
    .Q(\lfsr0.stop_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3028_ (.CLK(clknet_leaf_20_clk),
    .D(net418),
    .RESET_B(net79),
    .Q(\lfsr0.stop_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3029_ (.CLK(clknet_leaf_19_clk),
    .D(_0357_),
    .RESET_B(net91),
    .Q(\lfsr0.stop_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3030_ (.CLK(clknet_leaf_2_clk),
    .D(net395),
    .RESET_B(net85),
    .Q(\lfsr0.stop_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3031_ (.CLK(clknet_leaf_1_clk),
    .D(_0359_),
    .RESET_B(net85),
    .Q(\lfsr0.stop_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3032_ (.CLK(clknet_leaf_2_clk),
    .D(net451),
    .RESET_B(net98),
    .Q(\lfsr0.stop_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3033_ (.CLK(clknet_leaf_3_clk),
    .D(_0361_),
    .RESET_B(net97),
    .Q(\lfsr0.stop_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3034_ (.CLK(clknet_leaf_3_clk),
    .D(_0362_),
    .RESET_B(net96),
    .Q(\lfsr0.stop_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3035_ (.CLK(clknet_leaf_2_clk),
    .D(_0363_),
    .RESET_B(net98),
    .Q(\lfsr0.stop_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3036_ (.CLK(clknet_leaf_1_clk),
    .D(_0364_),
    .RESET_B(net83),
    .Q(\lfsr0.stop_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3037_ (.CLK(clknet_leaf_20_clk),
    .D(_0365_),
    .RESET_B(net84),
    .Q(\lfsr0.stop_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _3038_ (.CLK(clknet_leaf_23_clk),
    .D(_0366_),
    .RESET_B(net80),
    .Q(\lfsr0.stop_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _3039_ (.CLK(clknet_leaf_23_clk),
    .D(net421),
    .RESET_B(net81),
    .Q(\lfsr0.stop_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _3040_ (.CLK(clknet_leaf_23_clk),
    .D(_0368_),
    .RESET_B(net80),
    .Q(\lfsr0.stop_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _3041_ (.CLK(clknet_leaf_0_clk),
    .D(_0369_),
    .RESET_B(net81),
    .Q(\lfsr0.stop_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _3042_ (.CLK(clknet_leaf_3_clk),
    .D(_0370_),
    .RESET_B(net97),
    .Q(\lfsr0.stop_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _3043_ (.CLK(clknet_leaf_3_clk),
    .D(_0371_),
    .RESET_B(net95),
    .Q(\lfsr0.stop_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _3044_ (.CLK(clknet_leaf_4_clk),
    .D(_0372_),
    .RESET_B(net94),
    .Q(\lfsr0.stop_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _3045_ (.CLK(clknet_leaf_4_clk),
    .D(_0373_),
    .RESET_B(net93),
    .Q(\lfsr0.stop_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _3046_ (.CLK(clknet_leaf_0_clk),
    .D(net425),
    .RESET_B(net93),
    .Q(\lfsr0.stop_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _3047_ (.CLK(clknet_leaf_0_clk),
    .D(_0375_),
    .RESET_B(net82),
    .Q(\lfsr0.stop_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _3048_ (.CLK(clknet_leaf_0_clk),
    .D(net415),
    .RESET_B(net81),
    .Q(\lfsr0.stop_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _3049_ (.CLK(clknet_leaf_0_clk),
    .D(net427),
    .RESET_B(net82),
    .Q(\lfsr0.stop_reg[23] ));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_138 (.HI(net138));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_139 (.HI(net139));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_140 (.HI(net140));
 sky130_fd_sc_hd__inv_2 _1376__1 (.A(clknet_2_2__leaf_ui_in[1]),
    .Y(net141));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 _2705__137 (.HI(net137));
 sky130_fd_sc_hd__buf_2 _3067_ (.A(\gray_sobel0.select_sobel_mux ),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _3068_ (.A(net76),
    .X(uo_out[1]));
 sky130_fd_sc_hd__clkbuf_4 _3069_ (.A(net200),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _3070_ (.A(\spi0.spi0.sdo_o ),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _3071_ (.A(\lfsr0.lfsr_done ),
    .X(uo_out[4]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(net171),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(net192),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(net194),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net180),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net188),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(net196),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net178),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net184),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(net174),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(net182),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(net190),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(net176),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net186),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net16),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(_0387_),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net19),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(_0386_),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net22),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(_0380_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(_1002_),
    .X(net23));
 sky130_fd_sc_hd__buf_1 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(_1002_),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(_0001_),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net32),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(_1211_),
    .X(net32));
 sky130_fd_sc_hd__buf_4 fanout33 (.A(\gray_sobel0.sobel0.next[0] ),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(_0485_),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout36 (.A(_0485_),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(_0484_),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout39 (.A(_0484_),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(_0433_),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(_0433_),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net45),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(\gray_sobel0.sobel0.next[1] ),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net49),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout49 (.A(\gray_sobel0.sobel0.next[1] ),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net53),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net53),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(_0008_),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__buf_4 fanout55 (.A(_1138_),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(_1138_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net59),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(_1139_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net62),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(_0384_),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(net65),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(\spi0.rxtx_done_rising ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net68),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(\lfsr0.lfsr_en_i ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(net71),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(\lfsr0.config_i ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net75),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(LFSR_enable_i_sync),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(\sgnl_sync1.signal_o ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(\gray_sobel0.select_sobel_mux ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net80),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net92),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(net83),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(net92),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(net92),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net92),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(net88),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(net91),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(net114),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 fanout93 (.A(net96),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 fanout94 (.A(net96),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout96 (.A(net99),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 fanout97 (.A(net99),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(net114),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 fanout101 (.A(net114),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(net114),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_2 fanout106 (.A(net113),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net113),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(net113),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net112),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_2 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net246),
    .X(net114));
 sky130_fd_sc_hd__buf_4 fanout115 (.A(net117),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(net193),
    .X(net117));
 sky130_fd_sc_hd__buf_4 fanout118 (.A(net121),
    .X(net118));
 sky130_fd_sc_hd__buf_2 fanout119 (.A(net121),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(net193),
    .X(net123));
 sky130_fd_sc_hd__conb_1 tt_um_gray_sobel_124 (.LO(net124));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__bufinv_16 clkload3 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload5 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__inv_8 clkload8 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__inv_12 clkload9 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload10 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__inv_12 clkload11 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload12 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__inv_12 clkload14 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__inv_8 clkload15 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkinv_8 clkload16 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinv_4 clkload17 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_4 clkload18 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__inv_8 clkload19 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__inv_6 clkload20 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__inv_6 clkload21 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__inv_12 clkload22 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_ui_in[1]  (.A(ui_in[1]),
    .X(clknet_0_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_2_0__leaf_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_2_1__leaf_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_2_2__leaf_ui_in[1]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_ui_in[1]  (.A(clknet_0_ui_in[1]),
    .X(clknet_2_3__leaf_ui_in[1]));
 sky130_fd_sc_hd__clkinv_16 clkload23 (.A(clknet_2_0__leaf_ui_in[1]));
 sky130_fd_sc_hd__clkinv_16 clkload24 (.A(clknet_2_1__leaf_ui_in[1]));
 sky130_fd_sc_hd__inv_12 clkload25 (.A(clknet_2_3__leaf_ui_in[1]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net1),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(rst_n),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(uio_in[0]),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net9),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(uio_in[3]),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net12),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(ui_in[6]),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net7),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(ui_in[3]),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net4),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(uio_in[1]),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net10),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(ui_in[7]),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net8),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(uio_in[4]),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net13),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(ui_in[4]),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net5),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(uio_in[2]),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net11),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(ui_in[0]),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net2),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(ui_in[2]),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net3),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(ui_in[5]),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net6),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[5] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i2[3] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(ena),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[2] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[4] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[6] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[6] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\spi0.signal_sync1.signal_sync ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\nreset_sync0.r_sync ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\sgnl_sync3.signal_sync ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\sgnl_sync1.signal_sync ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\sgnl_sync8.signal_sync ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\sgnl_sync6.signal_sync ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\spi0.spi0.data_rx_o[1] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\sgnl_sync0.signal_sync ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\sgnl_sync4.signal_sync ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\sgnl_sync5.signal_sync ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\sgnl_sync7.signal_sync ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\sgnl_sync2.signal_sync ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\spi0.spi0.data_rx_o[21] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\spi0.spi0.data_rx_o[6] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\spi0.spi0.data_rx_o[18] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\spi0.spi0.data_rx_o[14] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\spi0.spi0.data_rx_o[13] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\spi0.rxtx_done ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\spi0.spi0.data_rx_o[7] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\spi0.spi0.data_rx_o[22] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\spi0.spi0.data_rx_o[17] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\spi0.spi0.data_rx_o[12] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\spi0.spi0.data_rx_o[16] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\spi0.spi0.data_rx_o[3] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\spi0.spi0.data_rx_o[10] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\spi0.spi0.data_rx_o[4] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\spi0.spi0.data_rx_o[15] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\spi0.spi0.data_rx_o[8] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\spi0.spi0.data_rx_o[11] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[7] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\spi0.spi0.data_rx_o[9] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\spi0.spi0.data_rx_o[5] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[7] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\spi0.spi0.data_rx_o[19] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\spi0.spi0.data_rx_o[20] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[6] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[3] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\spi0.spi0.data_rx_o[2] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[3] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[2] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[0] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\gray_sobel0.gray_scale0.nreset_i ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i5[0] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[2] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i1[1] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\spi0.spi0.sdo_register[22] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\spi0.spi0.sdo_register[16] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\spi0.spi0.sdo_register[7] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\spi0.spi0.sdo_register[15] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\spi0.spi0.sdo_register[18] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\spi0.spi0.sdo_register[8] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\spi0.spi0.sdo_register[11] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\spi0.spi0.sdo_register[1] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\spi0.spi0.sdo_register[6] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\spi0.spi0.sdo_register[13] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\spi0.spi0.sdo_register[20] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\spi0.spi0.sdo_register[4] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\spi0.spi0.sdo_register[3] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\spi0.spi0.sdo_register[9] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\spi0.spi0.sdo_register[17] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\spi0.spi0.sdo_register[21] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\spi0.spi0.sdo_register[2] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\sa0.en_i ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\spi0.spi0.sdo_register[5] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\spi0.spi0.sdo_register[10] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\spi0.spi0.sdo_register[19] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\spi0.spi0.sdo_register[12] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\spi0.spi0.sdo_register[14] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\spi0.spi0.sdo_register[0] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(lfsr_mode_sel_i_sync),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\spi0.spi0.counter[5] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\spi0.spi0.counter[0] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\gray_sobel0.out_px_sobel[7] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\spi0.spi0.counter[3] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\spi0.spi0.data_rx_o[0] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\spi0.data_tx[16] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[1] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\lfsr0.lfsr_rdy_o ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[2] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\gray_sobel0.out_px_sobel[0] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[4] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[5] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\spi0.data_tx[17] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[3] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\spi0.spi0.counter[2] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_1214_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[0] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\gray_sobel0.out_px_sobel[3] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[7] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\spi0.data_tx[7] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\spi0.data_tx[8] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\spi0.data_tx[23] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\gray_sobel0.sobel0.counter_pixels[23] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\spi0.data_tx[13] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\spi0.data_tx[15] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\spi0.data_tx[19] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\spi0.data_tx[22] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\spi0.data_tx[2] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\spi0.data_tx[5] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\spi0.data_tx[12] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\spi0.spi0.counter[1] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\spi0.data_tx[10] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\spi0.data_tx[0] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\spi0.data_tx[6] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\spi0.data_tx[3] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\spi0.data_tx[1] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\spi0.data_tx[4] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\spi0.data_tx[11] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\spi0.data_tx[21] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i4[6] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\gray_sobel0.out_px_sobel[1] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\spi0.data_tx[9] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\sa0.signature_o[23] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0197_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\gray_sobel0.out_px_sobel[4] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\lfsr0.seed_reg[15] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\lfsr0.seed_reg[10] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\lfsr0.seed_reg[20] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0350_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\lfsr0.seed_reg[1] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0331_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\gray_sobel0.out_px_sobel[5] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\lfsr0.seed_reg[0] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\lfsr0.seed_reg[6] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0336_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\spi0.data_tx[20] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\lfsr0.seed_reg[12] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\lfsr0.seed_reg[5] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0335_),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\spi0.data_tx[14] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\spi0.data_tx[18] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\lfsr0.seed_reg[13] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0343_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\gray_sobel0.out_px_sobel[6] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\lfsr0.seed_reg[18] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0348_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\lfsr0.seed_reg[17] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0347_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\lfsr0.seed_reg[9] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\lfsr0.seed_reg[22] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0352_),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\lfsr0.seed_reg[23] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0353_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\lfsr0.seed_reg[8] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\lfsr0.seed_reg[11] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\lfsr0.seed_reg[2] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0332_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\lfsr0.seed_reg[4] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_0334_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\lfsr0.seed_reg[14] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0344_),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\lfsr0.seed_reg[19] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0349_),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[6] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\sa0.signature_o[7] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\sa0.signature_o[17] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0192_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\lfsr0.seed_reg[21] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0351_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[7] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\sa0.signature_o[8] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\gray_sobel0.out_px_sobel[2] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\lfsr0.seed_reg[7] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\lfsr0.seed_reg[16] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0346_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\sa0.signature_o[11] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0186_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\gray_sobel0.sobel0.counter_pixels[17] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\gray_sobel0.sobel0.px_ready ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\gray_sobel0.sobel0.counter_pixels[5] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\lfsr0.seed_reg[3] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0333_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\sa0.signature_o[14] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0189_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\gray_sobel0.sobel0.counter_pixels[14] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\sa0.signature_o[15] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0190_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\sa0.signature_o[18] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0193_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\sa0.signature_o[16] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\sa0.signature_o[10] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\sa0.signature_o[19] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0194_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\sa0.signature_o[21] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0196_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\gray_sobel0.sobel0.counter_pixels[3] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[3] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\sa0.signature_o[20] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[2] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\input_data[4] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0358_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\sa0.signature_o[9] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\lfsr0.stop_reg[1] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0355_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\gray_sobel0.sobel0.counter_pixels[8] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\sa0.signature_o[12] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0187_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\gray_sobel0.sobel0.counter_pixels[20] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[7] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\sa0.signature_o[13] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\sa0.signature_o[6] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\sa0.signature_o[1] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\sa0.signature_o[3] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\gray_sobel0.sobel0.counter_pixels[6] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\sa0.signature_o[2] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\sa0.signature_o[5] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\input_data[3] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\input_data[16] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\sa0.signature_o[4] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\lfsr0.stop_reg[22] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0376_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[3] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\lfsr0.stop_reg[2] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0356_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i7[0] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\lfsr0.stop_reg[13] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0367_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\lfsr0.stop_reg[12] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\input_data[13] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\lfsr0.stop_reg[20] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0374_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\lfsr0.stop_reg[23] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0377_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\input_data[2] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\input_data[20] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i3[0] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\lfsr0.stop_reg[7] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\input_data[19] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\input_data[14] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\input_data[1] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\gray_sobel0.sobel0.counter_pixels[12] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\lfsr0.stop_reg[8] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\input_data[18] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i8[5] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\lfsr0.stop_reg[18] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(in_data_rdy),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\input_data[5] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\input_data[17] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\lfsr0.stop_reg[17] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\input_data[21] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\lfsr0.stop_reg[19] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\gray_sobel0.sobel0.counter_pixels[10] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\lfsr0.stop_reg[9] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\lfsr0.stop_reg[5] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\input_data[23] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\lfsr0.stop_reg[6] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0360_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\input_data[22] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\gray_sobel0.sobel0.sobel.matrix_pixels_i0[5] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\lfsr0.stop_reg[10] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\lfsr0.stop_reg[11] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\sa0.signature_o[0] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\lfsr0.stop_reg[15] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\input_data[6] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\gray_sobel0.sobel0.counter_pixels[9] ),
    .X(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\spi0.spi0.data_rx_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\spi0.spi0.data_rx_o[0] ));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_281 ();
 assign uio_oe[0] = net124;
 assign uio_oe[1] = net125;
 assign uio_oe[2] = net126;
 assign uio_oe[3] = net127;
 assign uio_oe[4] = net128;
 assign uio_oe[5] = net138;
 assign uio_oe[6] = net139;
 assign uio_oe[7] = net140;
 assign uio_out[0] = net129;
 assign uio_out[1] = net130;
 assign uio_out[2] = net131;
 assign uio_out[3] = net132;
 assign uio_out[4] = net133;
 assign uio_out[5] = net134;
 assign uio_out[6] = net135;
 assign uio_out[7] = net136;
endmodule
